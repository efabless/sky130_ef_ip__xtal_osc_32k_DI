VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_32k_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_32k_DI ;
  ORIGIN 0.000 0.000 ;
  SIZE 525.300 BY 211.800 ;
  PIN boost
    ANTENNAGATEAREA 0.510000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 219.330 75.500 219.500 76.000 ;
        RECT 220.300 75.500 220.470 76.000 ;
        RECT 220.355 71.080 220.685 71.570 ;
        RECT 215.825 67.310 215.995 67.640 ;
        RECT 217.420 67.310 217.590 67.640 ;
      LAYER mcon ;
        RECT 219.330 75.665 219.500 75.835 ;
        RECT 220.300 75.665 220.470 75.835 ;
        RECT 220.435 71.240 220.605 71.410 ;
        RECT 215.825 67.390 215.995 67.560 ;
        RECT 217.420 67.390 217.590 67.560 ;
      LAYER met1 ;
        RECT 217.390 75.820 217.720 75.870 ;
        RECT 219.300 75.820 219.530 75.980 ;
        RECT 220.270 75.820 220.500 75.980 ;
        RECT 217.390 75.620 220.500 75.820 ;
        RECT 217.390 75.280 217.720 75.620 ;
        RECT 219.290 75.520 219.530 75.620 ;
        RECT 220.270 75.520 220.500 75.620 ;
        RECT 217.475 71.480 217.745 71.845 ;
        RECT 220.325 71.480 220.715 71.550 ;
        RECT 217.475 71.220 220.715 71.480 ;
        RECT 217.475 71.170 217.745 71.220 ;
        RECT 220.325 71.100 220.715 71.220 ;
        RECT 215.795 67.550 216.025 67.620 ;
        RECT 216.440 67.550 216.810 67.600 ;
        RECT 217.390 67.550 217.620 67.620 ;
        RECT 215.780 67.310 217.640 67.550 ;
        RECT 216.440 67.130 216.810 67.310 ;
        RECT 216.130 66.130 217.130 67.130 ;
      LAYER via ;
        RECT 217.425 75.445 217.685 75.705 ;
        RECT 217.480 71.380 217.740 71.640 ;
        RECT 216.495 67.220 216.755 67.480 ;
      LAYER met2 ;
        RECT 217.340 75.330 217.770 75.820 ;
        RECT 217.430 71.795 217.700 75.330 ;
        RECT 217.425 71.220 217.795 71.795 ;
        RECT 217.430 68.490 217.700 71.220 ;
        RECT 216.495 68.220 217.700 68.490 ;
        RECT 216.495 67.865 216.765 68.220 ;
        RECT 216.495 67.550 216.810 67.865 ;
        RECT 216.390 67.150 216.860 67.550 ;
        RECT 216.540 64.930 216.810 67.150 ;
        RECT 216.195 0.000 217.195 64.930 ;
        RECT 216.195 -3.280 216.475 0.000 ;
    END
  END boost
  PIN ena
    ANTENNAGATEAREA 0.585000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 201.110 75.500 201.280 76.000 ;
        RECT 202.080 75.500 202.250 76.000 ;
        RECT 203.990 67.310 204.160 67.640 ;
        RECT 205.585 67.310 205.755 67.640 ;
        RECT 202.980 64.930 203.310 65.420 ;
        RECT 209.655 64.820 209.825 65.150 ;
      LAYER mcon ;
        RECT 201.110 75.665 201.280 75.835 ;
        RECT 202.080 75.665 202.250 75.835 ;
        RECT 203.990 67.390 204.160 67.560 ;
        RECT 205.585 67.390 205.755 67.560 ;
        RECT 203.060 65.090 203.230 65.260 ;
        RECT 209.655 64.900 209.825 65.070 ;
      LAYER met1 ;
        RECT 201.080 75.820 201.310 75.980 ;
        RECT 202.050 75.820 202.280 75.980 ;
        RECT 203.860 75.820 204.190 75.870 ;
        RECT 201.080 75.620 204.190 75.820 ;
        RECT 201.080 75.520 201.310 75.620 ;
        RECT 202.050 75.520 202.290 75.620 ;
        RECT 203.860 75.280 204.190 75.620 ;
        RECT 203.960 67.550 204.190 67.620 ;
        RECT 204.770 67.550 205.140 67.600 ;
        RECT 205.555 67.550 205.785 67.620 ;
        RECT 203.940 67.310 205.800 67.550 ;
        RECT 204.770 67.130 205.140 67.310 ;
        RECT 204.450 66.130 205.450 67.130 ;
        RECT 204.450 66.120 204.735 66.130 ;
        RECT 203.060 65.875 204.735 66.120 ;
        RECT 203.060 65.400 203.305 65.875 ;
        RECT 204.450 65.800 204.735 65.875 ;
        RECT 209.570 65.790 209.830 66.150 ;
        RECT 202.950 64.950 203.340 65.400 ;
        RECT 209.630 65.130 209.830 65.790 ;
        RECT 209.625 64.840 209.855 65.130 ;
      LAYER via ;
        RECT 203.895 75.445 204.155 75.705 ;
        RECT 204.825 67.220 205.085 67.480 ;
        RECT 204.465 65.875 204.725 66.135 ;
        RECT 209.570 65.840 209.830 66.100 ;
      LAYER met2 ;
        RECT 203.810 75.330 204.240 75.820 ;
        RECT 203.880 68.490 204.150 75.330 ;
        RECT 203.880 68.220 205.085 68.490 ;
        RECT 204.815 67.550 205.085 68.220 ;
        RECT 204.720 67.150 205.190 67.550 ;
        RECT 204.400 66.100 204.785 66.150 ;
        RECT 204.400 65.905 209.920 66.100 ;
        RECT 204.400 65.855 204.785 65.905 ;
        RECT 204.450 64.930 204.735 65.855 ;
        RECT 209.520 65.840 209.880 65.905 ;
        RECT 203.780 0.000 204.780 64.930 ;
        RECT 203.780 -3.280 204.060 0.000 ;
    END
  END ena
  PIN out
    PORT
      LAYER li1 ;
        RECT 220.165 130.060 222.325 130.750 ;
      LAYER mcon ;
        RECT 220.260 130.140 222.230 130.670 ;
      LAYER met1 ;
        RECT 221.020 133.100 222.020 134.100 ;
        RECT 221.235 130.700 221.770 133.100 ;
        RECT 220.190 130.110 222.295 130.700 ;
      LAYER via ;
        RECT 221.225 133.325 221.805 133.905 ;
      LAYER met2 ;
        RECT 515.825 166.965 516.465 218.525 ;
        RECT 221.020 165.865 516.465 166.965 ;
        RECT 221.020 133.100 222.020 165.865 ;
    END
  END out
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER li1 ;
        RECT 211.885 90.280 212.055 90.780 ;
        RECT 218.545 90.040 219.005 90.210 ;
        RECT 208.610 88.900 208.780 89.400 ;
        RECT 199.550 88.055 199.880 88.545 ;
        RECT 147.105 84.500 149.265 84.850 ;
        RECT 199.535 84.785 199.865 85.275 ;
      LAYER mcon ;
        RECT 211.885 90.445 212.055 90.615 ;
        RECT 218.690 90.040 218.860 90.210 ;
        RECT 208.610 89.065 208.780 89.235 ;
        RECT 199.630 88.215 199.800 88.385 ;
        RECT 199.615 84.945 199.785 85.115 ;
        RECT 147.205 84.590 147.375 84.760 ;
        RECT 147.565 84.590 147.735 84.760 ;
        RECT 147.925 84.590 148.095 84.760 ;
        RECT 148.285 84.590 148.455 84.760 ;
        RECT 148.645 84.590 148.815 84.760 ;
        RECT 149.005 84.590 149.175 84.760 ;
      LAYER met1 ;
        RECT 145.170 133.100 146.170 134.100 ;
        RECT 145.425 83.415 145.860 133.100 ;
        RECT 211.855 90.590 212.085 90.760 ;
        RECT 210.160 90.385 212.085 90.590 ;
        RECT 208.580 89.250 208.810 89.380 ;
        RECT 210.160 89.250 210.365 90.385 ;
        RECT 211.855 90.300 212.085 90.385 ;
        RECT 218.565 90.010 218.985 90.240 ;
        RECT 208.580 89.235 210.365 89.250 ;
        RECT 214.390 89.235 215.275 89.340 ;
        RECT 208.580 89.045 215.275 89.235 ;
        RECT 208.580 88.920 208.810 89.045 ;
        RECT 210.105 89.030 215.275 89.045 ;
        RECT 199.535 88.525 199.880 88.565 ;
        RECT 199.520 88.075 199.910 88.525 ;
        RECT 199.535 85.255 199.880 88.075 ;
        RECT 210.105 87.700 210.420 89.030 ;
        RECT 214.390 88.885 215.275 89.030 ;
        RECT 216.645 89.280 217.530 89.335 ;
        RECT 218.625 89.280 218.865 90.010 ;
        RECT 216.645 89.040 218.865 89.280 ;
        RECT 216.645 88.880 217.530 89.040 ;
        RECT 210.115 85.360 210.430 86.575 ;
        RECT 147.105 83.415 149.265 84.850 ;
        RECT 199.505 84.805 199.895 85.255 ;
        RECT 199.535 83.415 199.880 84.805 ;
        RECT 210.140 84.345 210.410 85.360 ;
        RECT 145.425 83.385 199.880 83.415 ;
        RECT 205.210 84.075 210.410 84.345 ;
        RECT 205.210 83.385 205.480 84.075 ;
        RECT 145.425 83.115 205.480 83.385 ;
        RECT 145.425 83.030 199.880 83.115 ;
        RECT 145.425 82.980 199.875 83.030 ;
      LAYER via ;
        RECT 145.385 133.325 145.965 133.905 ;
        RECT 214.545 88.985 214.805 89.245 ;
        RECT 214.865 88.985 215.125 89.245 ;
        RECT 216.800 88.980 217.060 89.240 ;
        RECT 217.120 88.980 217.380 89.240 ;
        RECT 210.135 88.500 210.395 88.760 ;
        RECT 210.135 88.180 210.395 88.440 ;
        RECT 210.135 87.860 210.395 88.120 ;
        RECT 210.145 86.160 210.405 86.420 ;
        RECT 210.145 85.840 210.405 86.100 ;
        RECT 210.145 85.520 210.405 85.780 ;
      LAYER met2 ;
        RECT 6.825 143.320 7.465 218.525 ;
        RECT 6.825 142.320 146.175 143.320 ;
        RECT 145.170 133.100 146.170 142.320 ;
        RECT 214.340 89.245 215.325 89.290 ;
        RECT 216.595 89.245 217.580 89.285 ;
        RECT 214.340 89.005 217.580 89.245 ;
        RECT 214.340 88.935 215.325 89.005 ;
        RECT 216.595 88.930 217.580 89.005 ;
        RECT 210.055 87.750 210.470 88.865 ;
        RECT 210.075 86.525 210.450 87.750 ;
        RECT 210.065 85.410 210.480 86.525 ;
    END
  END in
  PIN dout
    PORT
      LAYER li1 ;
        RECT 203.795 70.320 205.955 71.010 ;
      LAYER mcon ;
        RECT 203.890 70.400 205.860 70.930 ;
      LAYER met1 ;
        RECT 203.825 70.865 205.930 70.960 ;
        RECT 199.855 70.480 205.930 70.865 ;
        RECT 199.855 64.930 200.240 70.480 ;
        RECT 203.825 70.370 205.930 70.480 ;
        RECT 199.580 63.930 200.580 64.930 ;
      LAYER via ;
        RECT 199.775 64.155 200.355 64.735 ;
      LAYER met2 ;
        RECT 199.580 0.000 200.580 64.930 ;
        RECT 199.580 -3.280 199.860 0.000 ;
    END
  END dout
  PIN vdda1
    ANTENNADIFFAREA 200.228592 ;
    PORT
      LAYER nwell ;
        RECT 144.275 132.520 277.065 134.100 ;
        RECT 144.275 65.510 145.855 132.520 ;
        RECT 198.785 84.115 200.615 85.945 ;
        RECT 203.435 84.070 209.865 99.930 ;
        RECT 203.490 77.250 218.090 80.330 ;
        RECT 203.500 74.060 218.080 77.250 ;
        RECT 197.305 72.480 224.065 74.060 ;
        RECT 197.305 65.510 198.885 72.480 ;
        RECT 144.275 63.930 198.885 65.510 ;
        RECT 222.485 65.510 224.065 72.480 ;
        RECT 275.335 65.510 277.065 132.520 ;
        RECT 222.485 63.930 277.065 65.510 ;
      LAYER li1 ;
        RECT 151.175 133.665 171.595 133.815 ;
        RECT 172.625 133.665 192.445 133.770 ;
        RECT 193.180 133.665 219.810 133.815 ;
        RECT 249.865 133.665 269.770 133.765 ;
        RECT 271.995 133.665 274.145 133.770 ;
        RECT 144.710 133.495 276.630 133.665 ;
        RECT 144.710 130.945 144.880 133.495 ;
        RECT 151.175 133.395 171.595 133.495 ;
        RECT 172.625 133.395 192.445 133.495 ;
        RECT 193.180 133.380 219.810 133.495 ;
        RECT 249.865 133.390 269.770 133.495 ;
        RECT 271.995 133.395 274.145 133.495 ;
        RECT 276.460 133.225 276.630 133.495 ;
        RECT 271.995 131.200 274.155 131.550 ;
        RECT 144.605 65.265 144.935 130.945 ;
        RECT 209.365 99.540 209.970 99.560 ;
        RECT 207.215 99.505 209.970 99.540 ;
        RECT 203.020 99.370 209.970 99.505 ;
        RECT 203.020 97.410 207.385 99.370 ;
        RECT 209.305 97.410 209.970 99.370 ;
        RECT 203.020 96.290 209.970 97.410 ;
        RECT 203.020 94.330 203.995 96.290 ;
        RECT 204.905 95.620 205.365 95.790 ;
        RECT 205.915 94.330 207.385 96.290 ;
        RECT 209.305 94.330 209.970 96.290 ;
        RECT 203.020 93.210 209.970 94.330 ;
        RECT 203.020 91.250 203.995 93.210 ;
        RECT 204.905 92.540 205.365 92.710 ;
        RECT 205.915 91.250 207.385 93.210 ;
        RECT 209.305 91.250 209.970 93.210 ;
        RECT 203.020 90.130 209.970 91.250 ;
        RECT 203.020 88.170 203.995 90.130 ;
        RECT 204.905 89.460 205.365 89.630 ;
        RECT 205.915 88.170 207.385 90.130 ;
        RECT 209.305 88.170 209.970 90.130 ;
        RECT 203.020 87.050 209.970 88.170 ;
        RECT 198.965 85.760 200.435 85.765 ;
        RECT 198.965 85.595 200.675 85.760 ;
        RECT 198.965 84.465 199.135 85.595 ;
        RECT 200.265 84.465 200.675 85.595 ;
        RECT 198.965 84.295 200.675 84.465 ;
        RECT 203.020 85.090 203.995 87.050 ;
        RECT 204.905 85.590 205.365 85.760 ;
        RECT 205.915 85.090 207.385 87.050 ;
        RECT 207.935 85.590 208.395 85.760 ;
        RECT 209.305 85.090 209.970 87.050 ;
        RECT 203.020 84.420 209.970 85.090 ;
        RECT 200.265 84.290 200.675 84.295 ;
        RECT 203.530 79.730 210.280 80.360 ;
        RECT 203.530 77.810 204.070 79.730 ;
        RECT 206.320 77.810 207.400 79.730 ;
        RECT 208.305 78.310 208.765 78.480 ;
        RECT 209.660 77.810 210.280 79.730 ;
        RECT 203.530 76.720 210.280 77.810 ;
        RECT 203.530 74.760 204.070 76.720 ;
        RECT 206.330 76.690 210.280 76.720 ;
        RECT 206.330 74.760 207.400 76.690 ;
        RECT 208.305 76.020 208.765 76.190 ;
        RECT 203.530 74.750 207.400 74.760 ;
        RECT 209.660 74.750 210.280 76.690 ;
        RECT 203.530 74.120 210.280 74.750 ;
        RECT 211.300 79.730 218.050 80.360 ;
        RECT 211.300 77.810 211.920 79.730 ;
        RECT 212.815 78.310 213.275 78.480 ;
        RECT 214.180 77.810 215.260 79.730 ;
        RECT 217.510 77.810 218.050 79.730 ;
        RECT 211.300 76.720 218.050 77.810 ;
        RECT 211.300 76.690 215.250 76.720 ;
        RECT 211.300 74.750 211.920 76.690 ;
        RECT 212.815 76.020 213.275 76.190 ;
        RECT 214.180 74.760 215.250 76.690 ;
        RECT 217.510 74.760 218.050 76.720 ;
        RECT 214.180 74.750 218.050 74.760 ;
        RECT 211.300 74.120 218.050 74.750 ;
        RECT 198.710 73.135 222.745 73.200 ;
        RECT 198.270 72.965 223.150 73.135 ;
        RECT 198.270 72.235 198.440 72.965 ;
        RECT 198.710 72.900 222.745 72.965 ;
        RECT 222.980 72.395 223.150 72.965 ;
        RECT 147.155 66.560 149.315 66.910 ;
        RECT 144.710 64.535 144.880 65.265 ;
        RECT 198.185 64.905 198.505 72.235 ;
        RECT 222.885 65.210 223.175 72.395 ;
        RECT 147.155 64.535 149.310 64.640 ;
        RECT 151.135 64.535 171.045 64.625 ;
        RECT 172.645 64.535 192.475 64.635 ;
        RECT 193.225 64.535 197.880 64.645 ;
        RECT 198.270 64.535 198.440 64.905 ;
        RECT 144.710 64.365 198.440 64.535 ;
        RECT 222.980 64.535 223.150 65.210 ;
        RECT 276.345 64.835 276.725 133.225 ;
        RECT 223.850 64.535 248.185 64.665 ;
        RECT 249.925 64.535 269.755 64.630 ;
        RECT 276.460 64.535 276.630 64.835 ;
        RECT 222.980 64.365 276.630 64.535 ;
        RECT 147.155 64.265 149.310 64.365 ;
        RECT 151.135 64.255 171.045 64.365 ;
        RECT 172.645 64.265 192.475 64.365 ;
        RECT 193.225 64.270 197.880 64.365 ;
        RECT 223.850 64.350 248.185 64.365 ;
        RECT 249.925 64.265 269.755 64.365 ;
      LAYER mcon ;
        RECT 151.220 133.520 151.390 133.690 ;
        RECT 151.580 133.520 151.750 133.690 ;
        RECT 151.940 133.520 152.110 133.690 ;
        RECT 152.300 133.520 152.470 133.690 ;
        RECT 152.660 133.520 152.830 133.690 ;
        RECT 153.020 133.520 153.190 133.690 ;
        RECT 153.380 133.520 153.550 133.690 ;
        RECT 153.740 133.520 153.910 133.690 ;
        RECT 154.100 133.520 154.270 133.690 ;
        RECT 154.460 133.520 154.630 133.690 ;
        RECT 154.820 133.520 154.990 133.690 ;
        RECT 155.180 133.520 155.350 133.690 ;
        RECT 155.540 133.520 155.710 133.690 ;
        RECT 155.900 133.520 156.070 133.690 ;
        RECT 156.260 133.520 156.430 133.690 ;
        RECT 156.620 133.520 156.790 133.690 ;
        RECT 156.980 133.520 157.150 133.690 ;
        RECT 157.340 133.520 157.510 133.690 ;
        RECT 157.700 133.520 157.870 133.690 ;
        RECT 158.060 133.520 158.230 133.690 ;
        RECT 158.420 133.520 158.590 133.690 ;
        RECT 158.780 133.520 158.950 133.690 ;
        RECT 159.140 133.520 159.310 133.690 ;
        RECT 159.500 133.520 159.670 133.690 ;
        RECT 159.860 133.520 160.030 133.690 ;
        RECT 160.220 133.520 160.390 133.690 ;
        RECT 160.580 133.520 160.750 133.690 ;
        RECT 160.940 133.520 161.110 133.690 ;
        RECT 161.300 133.520 161.470 133.690 ;
        RECT 161.660 133.520 161.830 133.690 ;
        RECT 162.020 133.520 162.190 133.690 ;
        RECT 162.380 133.520 162.550 133.690 ;
        RECT 162.740 133.520 162.910 133.690 ;
        RECT 163.100 133.520 163.270 133.690 ;
        RECT 163.460 133.520 163.630 133.690 ;
        RECT 163.820 133.520 163.990 133.690 ;
        RECT 164.180 133.520 164.350 133.690 ;
        RECT 164.540 133.520 164.710 133.690 ;
        RECT 164.900 133.520 165.070 133.690 ;
        RECT 165.260 133.520 165.430 133.690 ;
        RECT 165.620 133.520 165.790 133.690 ;
        RECT 165.980 133.520 166.150 133.690 ;
        RECT 166.340 133.520 166.510 133.690 ;
        RECT 166.700 133.520 166.870 133.690 ;
        RECT 167.060 133.520 167.230 133.690 ;
        RECT 167.420 133.520 167.590 133.690 ;
        RECT 167.780 133.520 167.950 133.690 ;
        RECT 168.140 133.520 168.310 133.690 ;
        RECT 168.500 133.520 168.670 133.690 ;
        RECT 168.860 133.520 169.030 133.690 ;
        RECT 169.220 133.520 169.390 133.690 ;
        RECT 169.580 133.520 169.750 133.690 ;
        RECT 169.940 133.520 170.110 133.690 ;
        RECT 170.300 133.520 170.470 133.690 ;
        RECT 170.660 133.520 170.830 133.690 ;
        RECT 171.020 133.520 171.190 133.690 ;
        RECT 171.380 133.520 171.550 133.690 ;
        RECT 172.730 133.500 172.900 133.670 ;
        RECT 173.090 133.500 173.260 133.670 ;
        RECT 173.450 133.500 173.620 133.670 ;
        RECT 173.810 133.500 173.980 133.670 ;
        RECT 174.170 133.500 174.340 133.670 ;
        RECT 174.530 133.500 174.700 133.670 ;
        RECT 174.890 133.500 175.060 133.670 ;
        RECT 175.250 133.500 175.420 133.670 ;
        RECT 175.610 133.500 175.780 133.670 ;
        RECT 175.970 133.500 176.140 133.670 ;
        RECT 176.330 133.500 176.500 133.670 ;
        RECT 176.690 133.500 176.860 133.670 ;
        RECT 177.050 133.500 177.220 133.670 ;
        RECT 177.410 133.500 177.580 133.670 ;
        RECT 177.770 133.500 177.940 133.670 ;
        RECT 178.130 133.500 178.300 133.670 ;
        RECT 178.490 133.500 178.660 133.670 ;
        RECT 178.850 133.500 179.020 133.670 ;
        RECT 179.210 133.500 179.380 133.670 ;
        RECT 179.570 133.500 179.740 133.670 ;
        RECT 179.930 133.500 180.100 133.670 ;
        RECT 180.290 133.500 180.460 133.670 ;
        RECT 180.650 133.500 180.820 133.670 ;
        RECT 181.010 133.500 181.180 133.670 ;
        RECT 181.370 133.500 181.540 133.670 ;
        RECT 181.730 133.500 181.900 133.670 ;
        RECT 182.090 133.500 182.260 133.670 ;
        RECT 182.450 133.500 182.620 133.670 ;
        RECT 182.810 133.500 182.980 133.670 ;
        RECT 183.170 133.500 183.340 133.670 ;
        RECT 183.530 133.500 183.700 133.670 ;
        RECT 183.890 133.500 184.060 133.670 ;
        RECT 184.250 133.500 184.420 133.670 ;
        RECT 184.610 133.500 184.780 133.670 ;
        RECT 184.970 133.500 185.140 133.670 ;
        RECT 185.330 133.500 185.500 133.670 ;
        RECT 185.690 133.500 185.860 133.670 ;
        RECT 186.050 133.500 186.220 133.670 ;
        RECT 186.410 133.500 186.580 133.670 ;
        RECT 186.770 133.500 186.940 133.670 ;
        RECT 187.130 133.500 187.300 133.670 ;
        RECT 187.490 133.500 187.660 133.670 ;
        RECT 187.850 133.500 188.020 133.670 ;
        RECT 188.210 133.500 188.380 133.670 ;
        RECT 188.570 133.500 188.740 133.670 ;
        RECT 188.930 133.500 189.100 133.670 ;
        RECT 189.290 133.500 189.460 133.670 ;
        RECT 189.650 133.500 189.820 133.670 ;
        RECT 190.010 133.500 190.180 133.670 ;
        RECT 190.370 133.500 190.540 133.670 ;
        RECT 190.730 133.500 190.900 133.670 ;
        RECT 191.090 133.500 191.260 133.670 ;
        RECT 191.450 133.500 191.620 133.670 ;
        RECT 191.810 133.500 191.980 133.670 ;
        RECT 192.170 133.500 192.340 133.670 ;
        RECT 193.270 133.515 193.440 133.685 ;
        RECT 193.630 133.515 193.800 133.685 ;
        RECT 193.990 133.515 194.160 133.685 ;
        RECT 194.350 133.515 194.520 133.685 ;
        RECT 194.710 133.515 194.880 133.685 ;
        RECT 195.070 133.515 195.240 133.685 ;
        RECT 195.430 133.515 195.600 133.685 ;
        RECT 195.790 133.515 195.960 133.685 ;
        RECT 196.150 133.515 196.320 133.685 ;
        RECT 196.510 133.515 196.680 133.685 ;
        RECT 196.870 133.515 197.040 133.685 ;
        RECT 197.230 133.515 197.400 133.685 ;
        RECT 197.590 133.515 197.760 133.685 ;
        RECT 197.950 133.515 198.120 133.685 ;
        RECT 198.310 133.515 198.480 133.685 ;
        RECT 198.670 133.515 198.840 133.685 ;
        RECT 199.030 133.515 199.200 133.685 ;
        RECT 199.390 133.515 199.560 133.685 ;
        RECT 199.750 133.515 199.920 133.685 ;
        RECT 200.110 133.515 200.280 133.685 ;
        RECT 200.470 133.515 200.640 133.685 ;
        RECT 200.830 133.515 201.000 133.685 ;
        RECT 201.190 133.515 201.360 133.685 ;
        RECT 201.550 133.515 201.720 133.685 ;
        RECT 201.910 133.515 202.080 133.685 ;
        RECT 202.270 133.515 202.440 133.685 ;
        RECT 202.630 133.515 202.800 133.685 ;
        RECT 202.990 133.515 203.160 133.685 ;
        RECT 203.350 133.515 203.520 133.685 ;
        RECT 203.710 133.515 203.880 133.685 ;
        RECT 204.070 133.515 204.240 133.685 ;
        RECT 204.430 133.515 204.600 133.685 ;
        RECT 204.790 133.515 204.960 133.685 ;
        RECT 205.150 133.515 205.320 133.685 ;
        RECT 205.510 133.515 205.680 133.685 ;
        RECT 205.870 133.515 206.040 133.685 ;
        RECT 206.230 133.515 206.400 133.685 ;
        RECT 206.590 133.515 206.760 133.685 ;
        RECT 206.950 133.515 207.120 133.685 ;
        RECT 207.310 133.515 207.480 133.685 ;
        RECT 207.670 133.515 207.840 133.685 ;
        RECT 208.030 133.515 208.200 133.685 ;
        RECT 208.390 133.515 208.560 133.685 ;
        RECT 208.750 133.515 208.920 133.685 ;
        RECT 209.110 133.515 209.280 133.685 ;
        RECT 209.470 133.515 209.640 133.685 ;
        RECT 209.830 133.515 210.000 133.685 ;
        RECT 210.190 133.515 210.360 133.685 ;
        RECT 210.550 133.515 210.720 133.685 ;
        RECT 210.910 133.515 211.080 133.685 ;
        RECT 211.270 133.515 211.440 133.685 ;
        RECT 211.630 133.515 211.800 133.685 ;
        RECT 211.990 133.515 212.160 133.685 ;
        RECT 212.350 133.515 212.520 133.685 ;
        RECT 212.710 133.515 212.880 133.685 ;
        RECT 213.070 133.515 213.240 133.685 ;
        RECT 213.430 133.515 213.600 133.685 ;
        RECT 213.790 133.515 213.960 133.685 ;
        RECT 214.150 133.515 214.320 133.685 ;
        RECT 214.510 133.515 214.680 133.685 ;
        RECT 214.870 133.515 215.040 133.685 ;
        RECT 215.230 133.515 215.400 133.685 ;
        RECT 215.590 133.515 215.760 133.685 ;
        RECT 215.950 133.515 216.120 133.685 ;
        RECT 216.310 133.515 216.480 133.685 ;
        RECT 216.670 133.515 216.840 133.685 ;
        RECT 217.030 133.515 217.200 133.685 ;
        RECT 217.390 133.515 217.560 133.685 ;
        RECT 217.750 133.515 217.920 133.685 ;
        RECT 218.110 133.515 218.280 133.685 ;
        RECT 218.470 133.515 218.640 133.685 ;
        RECT 218.830 133.515 219.000 133.685 ;
        RECT 219.190 133.515 219.360 133.685 ;
        RECT 219.550 133.515 219.720 133.685 ;
        RECT 250.015 133.495 250.185 133.665 ;
        RECT 250.375 133.495 250.545 133.665 ;
        RECT 250.735 133.495 250.905 133.665 ;
        RECT 251.095 133.495 251.265 133.665 ;
        RECT 251.455 133.495 251.625 133.665 ;
        RECT 251.815 133.495 251.985 133.665 ;
        RECT 252.175 133.495 252.345 133.665 ;
        RECT 252.535 133.495 252.705 133.665 ;
        RECT 252.895 133.495 253.065 133.665 ;
        RECT 253.255 133.495 253.425 133.665 ;
        RECT 253.615 133.495 253.785 133.665 ;
        RECT 253.975 133.495 254.145 133.665 ;
        RECT 254.335 133.495 254.505 133.665 ;
        RECT 254.695 133.495 254.865 133.665 ;
        RECT 255.055 133.495 255.225 133.665 ;
        RECT 255.415 133.495 255.585 133.665 ;
        RECT 255.775 133.495 255.945 133.665 ;
        RECT 256.135 133.495 256.305 133.665 ;
        RECT 256.495 133.495 256.665 133.665 ;
        RECT 256.855 133.495 257.025 133.665 ;
        RECT 257.215 133.495 257.385 133.665 ;
        RECT 257.575 133.495 257.745 133.665 ;
        RECT 257.935 133.495 258.105 133.665 ;
        RECT 258.295 133.495 258.465 133.665 ;
        RECT 258.655 133.495 258.825 133.665 ;
        RECT 259.015 133.495 259.185 133.665 ;
        RECT 259.375 133.495 259.545 133.665 ;
        RECT 259.735 133.495 259.905 133.665 ;
        RECT 260.095 133.495 260.265 133.665 ;
        RECT 260.455 133.495 260.625 133.665 ;
        RECT 260.815 133.495 260.985 133.665 ;
        RECT 261.175 133.495 261.345 133.665 ;
        RECT 261.535 133.495 261.705 133.665 ;
        RECT 261.895 133.495 262.065 133.665 ;
        RECT 262.255 133.495 262.425 133.665 ;
        RECT 262.615 133.495 262.785 133.665 ;
        RECT 262.975 133.495 263.145 133.665 ;
        RECT 263.335 133.495 263.505 133.665 ;
        RECT 263.695 133.495 263.865 133.665 ;
        RECT 264.055 133.495 264.225 133.665 ;
        RECT 264.415 133.495 264.585 133.665 ;
        RECT 264.775 133.495 264.945 133.665 ;
        RECT 265.135 133.495 265.305 133.665 ;
        RECT 265.495 133.495 265.665 133.665 ;
        RECT 265.855 133.495 266.025 133.665 ;
        RECT 266.215 133.495 266.385 133.665 ;
        RECT 266.575 133.495 266.745 133.665 ;
        RECT 266.935 133.495 267.105 133.665 ;
        RECT 267.295 133.495 267.465 133.665 ;
        RECT 267.655 133.495 267.825 133.665 ;
        RECT 268.015 133.495 268.185 133.665 ;
        RECT 268.375 133.495 268.545 133.665 ;
        RECT 268.735 133.495 268.905 133.665 ;
        RECT 269.095 133.495 269.265 133.665 ;
        RECT 269.455 133.495 269.625 133.665 ;
        RECT 272.085 133.500 272.255 133.670 ;
        RECT 272.445 133.500 272.615 133.670 ;
        RECT 272.805 133.500 272.975 133.670 ;
        RECT 273.165 133.500 273.335 133.670 ;
        RECT 273.525 133.500 273.695 133.670 ;
        RECT 273.885 133.500 274.055 133.670 ;
        RECT 276.450 132.965 276.620 133.135 ;
        RECT 276.450 132.605 276.620 132.775 ;
        RECT 276.450 132.245 276.620 132.415 ;
        RECT 276.450 131.885 276.620 132.055 ;
        RECT 272.090 131.290 272.260 131.460 ;
        RECT 272.450 131.290 272.620 131.460 ;
        RECT 272.810 131.290 272.980 131.460 ;
        RECT 273.170 131.290 273.340 131.460 ;
        RECT 273.530 131.290 273.700 131.460 ;
        RECT 273.890 131.290 274.060 131.460 ;
        RECT 276.450 131.525 276.620 131.695 ;
        RECT 276.450 131.165 276.620 131.335 ;
        RECT 144.685 130.600 144.855 130.770 ;
        RECT 144.685 130.240 144.855 130.410 ;
        RECT 144.685 129.880 144.855 130.050 ;
        RECT 144.685 129.520 144.855 129.690 ;
        RECT 144.685 129.160 144.855 129.330 ;
        RECT 144.685 128.800 144.855 128.970 ;
        RECT 144.685 128.440 144.855 128.610 ;
        RECT 144.685 128.080 144.855 128.250 ;
        RECT 144.685 127.720 144.855 127.890 ;
        RECT 144.685 127.360 144.855 127.530 ;
        RECT 144.685 127.000 144.855 127.170 ;
        RECT 144.685 126.640 144.855 126.810 ;
        RECT 144.685 126.280 144.855 126.450 ;
        RECT 144.685 125.920 144.855 126.090 ;
        RECT 144.685 125.560 144.855 125.730 ;
        RECT 144.685 125.200 144.855 125.370 ;
        RECT 144.685 124.840 144.855 125.010 ;
        RECT 144.685 124.480 144.855 124.650 ;
        RECT 144.685 124.120 144.855 124.290 ;
        RECT 144.685 123.760 144.855 123.930 ;
        RECT 144.685 123.400 144.855 123.570 ;
        RECT 144.685 123.040 144.855 123.210 ;
        RECT 144.685 122.680 144.855 122.850 ;
        RECT 144.685 122.320 144.855 122.490 ;
        RECT 144.685 121.960 144.855 122.130 ;
        RECT 144.685 121.600 144.855 121.770 ;
        RECT 144.685 121.240 144.855 121.410 ;
        RECT 144.685 120.880 144.855 121.050 ;
        RECT 144.685 120.520 144.855 120.690 ;
        RECT 144.685 120.160 144.855 120.330 ;
        RECT 144.685 119.800 144.855 119.970 ;
        RECT 144.685 119.440 144.855 119.610 ;
        RECT 144.685 119.080 144.855 119.250 ;
        RECT 144.685 118.720 144.855 118.890 ;
        RECT 144.685 118.360 144.855 118.530 ;
        RECT 144.685 118.000 144.855 118.170 ;
        RECT 144.685 117.640 144.855 117.810 ;
        RECT 144.685 117.280 144.855 117.450 ;
        RECT 144.685 116.920 144.855 117.090 ;
        RECT 144.685 116.560 144.855 116.730 ;
        RECT 144.685 116.200 144.855 116.370 ;
        RECT 144.685 115.840 144.855 116.010 ;
        RECT 144.685 115.480 144.855 115.650 ;
        RECT 144.685 115.120 144.855 115.290 ;
        RECT 144.685 114.760 144.855 114.930 ;
        RECT 144.685 114.400 144.855 114.570 ;
        RECT 144.685 114.040 144.855 114.210 ;
        RECT 144.685 113.680 144.855 113.850 ;
        RECT 144.685 113.320 144.855 113.490 ;
        RECT 144.685 112.960 144.855 113.130 ;
        RECT 144.685 112.600 144.855 112.770 ;
        RECT 144.685 112.240 144.855 112.410 ;
        RECT 144.685 111.880 144.855 112.050 ;
        RECT 144.685 111.520 144.855 111.690 ;
        RECT 144.685 111.160 144.855 111.330 ;
        RECT 144.685 110.800 144.855 110.970 ;
        RECT 144.685 110.440 144.855 110.610 ;
        RECT 144.685 110.080 144.855 110.250 ;
        RECT 144.685 109.720 144.855 109.890 ;
        RECT 144.685 109.360 144.855 109.530 ;
        RECT 144.685 109.000 144.855 109.170 ;
        RECT 144.685 108.640 144.855 108.810 ;
        RECT 144.685 108.280 144.855 108.450 ;
        RECT 144.685 107.920 144.855 108.090 ;
        RECT 144.685 107.560 144.855 107.730 ;
        RECT 144.685 107.200 144.855 107.370 ;
        RECT 144.685 106.840 144.855 107.010 ;
        RECT 144.685 106.480 144.855 106.650 ;
        RECT 144.685 106.120 144.855 106.290 ;
        RECT 144.685 105.760 144.855 105.930 ;
        RECT 144.685 105.400 144.855 105.570 ;
        RECT 144.685 105.040 144.855 105.210 ;
        RECT 144.685 104.680 144.855 104.850 ;
        RECT 144.685 104.320 144.855 104.490 ;
        RECT 144.685 103.960 144.855 104.130 ;
        RECT 144.685 103.600 144.855 103.770 ;
        RECT 144.685 103.240 144.855 103.410 ;
        RECT 144.685 102.880 144.855 103.050 ;
        RECT 144.685 102.520 144.855 102.690 ;
        RECT 144.685 102.160 144.855 102.330 ;
        RECT 144.685 101.800 144.855 101.970 ;
        RECT 144.685 101.440 144.855 101.610 ;
        RECT 144.685 101.080 144.855 101.250 ;
        RECT 144.685 100.720 144.855 100.890 ;
        RECT 144.685 100.360 144.855 100.530 ;
        RECT 144.685 100.000 144.855 100.170 ;
        RECT 144.685 99.640 144.855 99.810 ;
        RECT 276.450 130.805 276.620 130.975 ;
        RECT 276.450 130.445 276.620 130.615 ;
        RECT 276.450 130.085 276.620 130.255 ;
        RECT 276.450 129.725 276.620 129.895 ;
        RECT 276.450 129.365 276.620 129.535 ;
        RECT 276.450 129.005 276.620 129.175 ;
        RECT 276.450 128.645 276.620 128.815 ;
        RECT 276.450 128.285 276.620 128.455 ;
        RECT 276.450 127.925 276.620 128.095 ;
        RECT 276.450 127.565 276.620 127.735 ;
        RECT 276.450 127.205 276.620 127.375 ;
        RECT 276.450 126.845 276.620 127.015 ;
        RECT 276.450 126.485 276.620 126.655 ;
        RECT 276.450 126.125 276.620 126.295 ;
        RECT 276.450 125.765 276.620 125.935 ;
        RECT 276.450 125.405 276.620 125.575 ;
        RECT 276.450 125.045 276.620 125.215 ;
        RECT 276.450 124.685 276.620 124.855 ;
        RECT 276.450 124.325 276.620 124.495 ;
        RECT 276.450 123.965 276.620 124.135 ;
        RECT 276.450 123.605 276.620 123.775 ;
        RECT 276.450 123.245 276.620 123.415 ;
        RECT 276.450 122.885 276.620 123.055 ;
        RECT 276.450 122.525 276.620 122.695 ;
        RECT 276.450 122.165 276.620 122.335 ;
        RECT 276.450 121.805 276.620 121.975 ;
        RECT 276.450 121.445 276.620 121.615 ;
        RECT 276.450 121.085 276.620 121.255 ;
        RECT 276.450 120.725 276.620 120.895 ;
        RECT 276.450 120.365 276.620 120.535 ;
        RECT 276.450 120.005 276.620 120.175 ;
        RECT 276.450 119.645 276.620 119.815 ;
        RECT 276.450 119.285 276.620 119.455 ;
        RECT 276.450 118.925 276.620 119.095 ;
        RECT 276.450 118.565 276.620 118.735 ;
        RECT 276.450 118.205 276.620 118.375 ;
        RECT 276.450 117.845 276.620 118.015 ;
        RECT 276.450 117.485 276.620 117.655 ;
        RECT 276.450 117.125 276.620 117.295 ;
        RECT 276.450 116.765 276.620 116.935 ;
        RECT 276.450 116.405 276.620 116.575 ;
        RECT 276.450 116.045 276.620 116.215 ;
        RECT 276.450 115.685 276.620 115.855 ;
        RECT 276.450 115.325 276.620 115.495 ;
        RECT 276.450 114.965 276.620 115.135 ;
        RECT 276.450 114.605 276.620 114.775 ;
        RECT 276.450 114.245 276.620 114.415 ;
        RECT 276.450 113.885 276.620 114.055 ;
        RECT 276.450 113.525 276.620 113.695 ;
        RECT 276.450 113.165 276.620 113.335 ;
        RECT 276.450 112.805 276.620 112.975 ;
        RECT 276.450 112.445 276.620 112.615 ;
        RECT 276.450 112.085 276.620 112.255 ;
        RECT 276.450 111.725 276.620 111.895 ;
        RECT 276.450 111.365 276.620 111.535 ;
        RECT 276.450 111.005 276.620 111.175 ;
        RECT 276.450 110.645 276.620 110.815 ;
        RECT 276.450 110.285 276.620 110.455 ;
        RECT 276.450 109.925 276.620 110.095 ;
        RECT 276.450 109.565 276.620 109.735 ;
        RECT 276.450 109.205 276.620 109.375 ;
        RECT 276.450 108.845 276.620 109.015 ;
        RECT 276.450 108.485 276.620 108.655 ;
        RECT 276.450 108.125 276.620 108.295 ;
        RECT 276.450 107.765 276.620 107.935 ;
        RECT 276.450 107.405 276.620 107.575 ;
        RECT 276.450 107.045 276.620 107.215 ;
        RECT 276.450 106.685 276.620 106.855 ;
        RECT 276.450 106.325 276.620 106.495 ;
        RECT 276.450 105.965 276.620 106.135 ;
        RECT 276.450 105.605 276.620 105.775 ;
        RECT 276.450 105.245 276.620 105.415 ;
        RECT 276.450 104.885 276.620 105.055 ;
        RECT 276.450 104.525 276.620 104.695 ;
        RECT 276.450 104.165 276.620 104.335 ;
        RECT 276.450 103.805 276.620 103.975 ;
        RECT 276.450 103.445 276.620 103.615 ;
        RECT 276.450 103.085 276.620 103.255 ;
        RECT 276.450 102.725 276.620 102.895 ;
        RECT 276.450 102.365 276.620 102.535 ;
        RECT 276.450 102.005 276.620 102.175 ;
        RECT 276.450 101.645 276.620 101.815 ;
        RECT 276.450 101.285 276.620 101.455 ;
        RECT 276.450 100.925 276.620 101.095 ;
        RECT 276.450 100.565 276.620 100.735 ;
        RECT 276.450 100.205 276.620 100.375 ;
        RECT 276.450 99.845 276.620 100.015 ;
        RECT 144.685 99.280 144.855 99.450 ;
        RECT 144.685 98.920 144.855 99.090 ;
        RECT 144.685 98.560 144.855 98.730 ;
        RECT 144.685 98.200 144.855 98.370 ;
        RECT 144.685 97.840 144.855 98.010 ;
        RECT 144.685 97.480 144.855 97.650 ;
        RECT 144.685 97.120 144.855 97.290 ;
        RECT 144.685 96.760 144.855 96.930 ;
        RECT 144.685 96.400 144.855 96.570 ;
        RECT 144.685 96.040 144.855 96.210 ;
        RECT 144.685 95.680 144.855 95.850 ;
        RECT 144.685 95.320 144.855 95.490 ;
        RECT 144.685 94.960 144.855 95.130 ;
        RECT 144.685 94.600 144.855 94.770 ;
        RECT 144.685 94.240 144.855 94.410 ;
        RECT 144.685 93.880 144.855 94.050 ;
        RECT 144.685 93.520 144.855 93.690 ;
        RECT 144.685 93.160 144.855 93.330 ;
        RECT 144.685 92.800 144.855 92.970 ;
        RECT 144.685 92.440 144.855 92.610 ;
        RECT 144.685 92.080 144.855 92.250 ;
        RECT 144.685 91.720 144.855 91.890 ;
        RECT 144.685 91.360 144.855 91.530 ;
        RECT 144.685 91.000 144.855 91.170 ;
        RECT 144.685 90.640 144.855 90.810 ;
        RECT 144.685 90.280 144.855 90.450 ;
        RECT 144.685 89.920 144.855 90.090 ;
        RECT 144.685 89.560 144.855 89.730 ;
        RECT 144.685 89.200 144.855 89.370 ;
        RECT 144.685 88.840 144.855 89.010 ;
        RECT 144.685 88.480 144.855 88.650 ;
        RECT 144.685 88.120 144.855 88.290 ;
        RECT 144.685 87.760 144.855 87.930 ;
        RECT 144.685 87.400 144.855 87.570 ;
        RECT 144.685 87.040 144.855 87.210 ;
        RECT 144.685 86.680 144.855 86.850 ;
        RECT 144.685 86.320 144.855 86.490 ;
        RECT 144.685 85.960 144.855 86.130 ;
        RECT 144.685 85.600 144.855 85.770 ;
        RECT 206.195 98.955 206.365 99.125 ;
        RECT 206.195 98.595 206.365 98.765 ;
        RECT 206.195 98.235 206.365 98.405 ;
        RECT 206.195 97.875 206.365 98.045 ;
        RECT 206.195 97.515 206.365 97.685 ;
        RECT 206.195 97.155 206.365 97.325 ;
        RECT 206.195 96.795 206.365 96.965 ;
        RECT 205.050 95.620 205.220 95.790 ;
        RECT 206.195 95.765 206.365 95.935 ;
        RECT 206.555 95.765 206.725 95.935 ;
        RECT 206.915 95.765 207.085 95.935 ;
        RECT 205.050 92.540 205.220 92.710 ;
        RECT 206.190 92.560 206.360 92.730 ;
        RECT 206.550 92.560 206.720 92.730 ;
        RECT 206.910 92.560 207.080 92.730 ;
        RECT 205.050 89.460 205.220 89.630 ;
        RECT 206.195 89.555 206.365 89.725 ;
        RECT 206.555 89.555 206.725 89.725 ;
        RECT 206.915 89.555 207.085 89.725 ;
        RECT 144.685 85.240 144.855 85.410 ;
        RECT 144.685 84.880 144.855 85.050 ;
        RECT 144.685 84.520 144.855 84.690 ;
        RECT 144.685 84.160 144.855 84.330 ;
        RECT 200.385 85.480 200.555 85.650 ;
        RECT 200.385 85.120 200.555 85.290 ;
        RECT 200.385 84.760 200.555 84.930 ;
        RECT 200.385 84.400 200.555 84.570 ;
        RECT 205.050 85.590 205.220 85.760 ;
        RECT 208.080 85.590 208.250 85.760 ;
        RECT 206.205 85.415 206.375 85.585 ;
        RECT 206.565 85.415 206.735 85.585 ;
        RECT 206.925 85.415 207.095 85.585 ;
        RECT 276.450 99.485 276.620 99.655 ;
        RECT 276.450 99.125 276.620 99.295 ;
        RECT 276.450 98.765 276.620 98.935 ;
        RECT 276.450 98.405 276.620 98.575 ;
        RECT 276.450 98.045 276.620 98.215 ;
        RECT 276.450 97.685 276.620 97.855 ;
        RECT 276.450 97.325 276.620 97.495 ;
        RECT 276.450 96.965 276.620 97.135 ;
        RECT 276.450 96.605 276.620 96.775 ;
        RECT 276.450 96.245 276.620 96.415 ;
        RECT 276.450 95.885 276.620 96.055 ;
        RECT 276.450 95.525 276.620 95.695 ;
        RECT 276.450 95.165 276.620 95.335 ;
        RECT 276.450 94.805 276.620 94.975 ;
        RECT 276.450 94.445 276.620 94.615 ;
        RECT 276.450 94.085 276.620 94.255 ;
        RECT 276.450 93.725 276.620 93.895 ;
        RECT 276.450 93.365 276.620 93.535 ;
        RECT 276.450 93.005 276.620 93.175 ;
        RECT 276.450 92.645 276.620 92.815 ;
        RECT 276.450 92.285 276.620 92.455 ;
        RECT 276.450 91.925 276.620 92.095 ;
        RECT 276.450 91.565 276.620 91.735 ;
        RECT 276.450 91.205 276.620 91.375 ;
        RECT 276.450 90.845 276.620 91.015 ;
        RECT 276.450 90.485 276.620 90.655 ;
        RECT 276.450 90.125 276.620 90.295 ;
        RECT 276.450 89.765 276.620 89.935 ;
        RECT 276.450 89.405 276.620 89.575 ;
        RECT 276.450 89.045 276.620 89.215 ;
        RECT 276.450 88.685 276.620 88.855 ;
        RECT 276.450 88.325 276.620 88.495 ;
        RECT 276.450 87.965 276.620 88.135 ;
        RECT 276.450 87.605 276.620 87.775 ;
        RECT 276.450 87.245 276.620 87.415 ;
        RECT 276.450 86.885 276.620 87.055 ;
        RECT 276.450 86.525 276.620 86.695 ;
        RECT 276.450 86.165 276.620 86.335 ;
        RECT 276.450 85.805 276.620 85.975 ;
        RECT 276.450 85.445 276.620 85.615 ;
        RECT 276.450 85.085 276.620 85.255 ;
        RECT 276.450 84.725 276.620 84.895 ;
        RECT 276.450 84.365 276.620 84.535 ;
        RECT 144.685 83.800 144.855 83.970 ;
        RECT 144.685 83.440 144.855 83.610 ;
        RECT 144.685 83.080 144.855 83.250 ;
        RECT 144.685 82.720 144.855 82.890 ;
        RECT 144.685 82.360 144.855 82.530 ;
        RECT 144.685 82.000 144.855 82.170 ;
        RECT 144.685 81.640 144.855 81.810 ;
        RECT 144.685 81.280 144.855 81.450 ;
        RECT 144.685 80.920 144.855 81.090 ;
        RECT 144.685 80.560 144.855 80.730 ;
        RECT 144.685 80.200 144.855 80.370 ;
        RECT 276.450 84.005 276.620 84.175 ;
        RECT 276.450 83.645 276.620 83.815 ;
        RECT 276.450 83.285 276.620 83.455 ;
        RECT 276.450 82.925 276.620 83.095 ;
        RECT 276.450 82.565 276.620 82.735 ;
        RECT 276.450 82.205 276.620 82.375 ;
        RECT 276.450 81.845 276.620 82.015 ;
        RECT 276.450 81.485 276.620 81.655 ;
        RECT 276.450 81.125 276.620 81.295 ;
        RECT 276.450 80.765 276.620 80.935 ;
        RECT 276.450 80.405 276.620 80.575 ;
        RECT 144.685 79.840 144.855 80.010 ;
        RECT 144.685 79.480 144.855 79.650 ;
        RECT 144.685 79.120 144.855 79.290 ;
        RECT 144.685 78.760 144.855 78.930 ;
        RECT 144.685 78.400 144.855 78.570 ;
        RECT 144.685 78.040 144.855 78.210 ;
        RECT 144.685 77.680 144.855 77.850 ;
        RECT 144.685 77.320 144.855 77.490 ;
        RECT 144.685 76.960 144.855 77.130 ;
        RECT 144.685 76.600 144.855 76.770 ;
        RECT 144.685 76.240 144.855 76.410 ;
        RECT 144.685 75.880 144.855 76.050 ;
        RECT 144.685 75.520 144.855 75.690 ;
        RECT 144.685 75.160 144.855 75.330 ;
        RECT 144.685 74.800 144.855 74.970 ;
        RECT 144.685 74.440 144.855 74.610 ;
        RECT 144.685 74.080 144.855 74.250 ;
        RECT 209.170 79.970 209.340 80.140 ;
        RECT 209.530 79.970 209.700 80.140 ;
        RECT 209.890 79.970 210.060 80.140 ;
        RECT 208.450 78.310 208.620 78.480 ;
        RECT 208.500 76.975 210.110 77.505 ;
        RECT 208.450 76.020 208.620 76.190 ;
        RECT 209.225 74.340 209.395 74.510 ;
        RECT 209.585 74.340 209.755 74.510 ;
        RECT 209.945 74.340 210.115 74.510 ;
        RECT 211.520 79.970 211.690 80.140 ;
        RECT 211.880 79.970 212.050 80.140 ;
        RECT 212.240 79.970 212.410 80.140 ;
        RECT 212.960 78.310 213.130 78.480 ;
        RECT 211.470 76.975 213.080 77.505 ;
        RECT 212.960 76.020 213.130 76.190 ;
        RECT 211.465 74.340 211.635 74.510 ;
        RECT 211.825 74.340 211.995 74.510 ;
        RECT 212.185 74.340 212.355 74.510 ;
        RECT 276.450 80.045 276.620 80.215 ;
        RECT 276.450 79.685 276.620 79.855 ;
        RECT 276.450 79.325 276.620 79.495 ;
        RECT 276.450 78.965 276.620 79.135 ;
        RECT 276.450 78.605 276.620 78.775 ;
        RECT 276.450 78.245 276.620 78.415 ;
        RECT 276.450 77.885 276.620 78.055 ;
        RECT 276.450 77.525 276.620 77.695 ;
        RECT 276.450 77.165 276.620 77.335 ;
        RECT 276.450 76.805 276.620 76.975 ;
        RECT 276.450 76.445 276.620 76.615 ;
        RECT 276.450 76.085 276.620 76.255 ;
        RECT 276.450 75.725 276.620 75.895 ;
        RECT 276.450 75.365 276.620 75.535 ;
        RECT 276.450 75.005 276.620 75.175 ;
        RECT 276.450 74.645 276.620 74.815 ;
        RECT 276.450 74.285 276.620 74.455 ;
        RECT 144.685 73.720 144.855 73.890 ;
        RECT 144.685 73.360 144.855 73.530 ;
        RECT 276.450 73.925 276.620 74.095 ;
        RECT 276.450 73.565 276.620 73.735 ;
        RECT 276.450 73.205 276.620 73.375 ;
        RECT 144.685 73.000 144.855 73.170 ;
        RECT 144.685 72.640 144.855 72.810 ;
        RECT 144.685 72.280 144.855 72.450 ;
        RECT 198.765 72.965 198.935 73.135 ;
        RECT 199.125 72.965 199.295 73.135 ;
        RECT 199.485 72.965 199.655 73.135 ;
        RECT 199.845 72.965 200.015 73.135 ;
        RECT 200.205 72.965 200.375 73.135 ;
        RECT 200.565 72.965 200.735 73.135 ;
        RECT 200.925 72.965 201.095 73.135 ;
        RECT 201.285 72.965 201.455 73.135 ;
        RECT 201.645 72.965 201.815 73.135 ;
        RECT 202.005 72.965 202.175 73.135 ;
        RECT 202.365 72.965 202.535 73.135 ;
        RECT 202.725 72.965 202.895 73.135 ;
        RECT 203.085 72.965 203.255 73.135 ;
        RECT 203.445 72.965 203.615 73.135 ;
        RECT 203.805 72.965 203.975 73.135 ;
        RECT 204.165 72.965 204.335 73.135 ;
        RECT 204.525 72.965 204.695 73.135 ;
        RECT 204.885 72.965 205.055 73.135 ;
        RECT 205.245 72.965 205.415 73.135 ;
        RECT 205.605 72.965 205.775 73.135 ;
        RECT 205.965 72.965 206.135 73.135 ;
        RECT 206.325 72.965 206.495 73.135 ;
        RECT 206.685 72.965 206.855 73.135 ;
        RECT 207.045 72.965 207.215 73.135 ;
        RECT 207.405 72.965 207.575 73.135 ;
        RECT 207.765 72.965 207.935 73.135 ;
        RECT 208.125 72.965 208.295 73.135 ;
        RECT 208.485 72.965 208.655 73.135 ;
        RECT 208.845 72.965 209.015 73.135 ;
        RECT 209.205 72.965 209.375 73.135 ;
        RECT 209.565 72.965 209.735 73.135 ;
        RECT 209.925 72.965 210.095 73.135 ;
        RECT 210.285 72.965 210.455 73.135 ;
        RECT 210.645 72.965 210.815 73.135 ;
        RECT 211.005 72.965 211.175 73.135 ;
        RECT 211.365 72.965 211.535 73.135 ;
        RECT 211.725 72.965 211.895 73.135 ;
        RECT 212.085 72.965 212.255 73.135 ;
        RECT 212.445 72.965 212.615 73.135 ;
        RECT 212.805 72.965 212.975 73.135 ;
        RECT 213.165 72.965 213.335 73.135 ;
        RECT 213.525 72.965 213.695 73.135 ;
        RECT 213.885 72.965 214.055 73.135 ;
        RECT 214.245 72.965 214.415 73.135 ;
        RECT 214.605 72.965 214.775 73.135 ;
        RECT 214.965 72.965 215.135 73.135 ;
        RECT 215.325 72.965 215.495 73.135 ;
        RECT 215.685 72.965 215.855 73.135 ;
        RECT 216.045 72.965 216.215 73.135 ;
        RECT 216.405 72.965 216.575 73.135 ;
        RECT 216.765 72.965 216.935 73.135 ;
        RECT 217.125 72.965 217.295 73.135 ;
        RECT 217.485 72.965 217.655 73.135 ;
        RECT 217.845 72.965 218.015 73.135 ;
        RECT 218.205 72.965 218.375 73.135 ;
        RECT 218.565 72.965 218.735 73.135 ;
        RECT 218.925 72.965 219.095 73.135 ;
        RECT 219.285 72.965 219.455 73.135 ;
        RECT 219.645 72.965 219.815 73.135 ;
        RECT 220.005 72.965 220.175 73.135 ;
        RECT 220.365 72.965 220.535 73.135 ;
        RECT 220.725 72.965 220.895 73.135 ;
        RECT 221.085 72.965 221.255 73.135 ;
        RECT 221.445 72.965 221.615 73.135 ;
        RECT 221.805 72.965 221.975 73.135 ;
        RECT 222.165 72.965 222.335 73.135 ;
        RECT 222.525 72.965 222.695 73.135 ;
        RECT 276.450 72.845 276.620 73.015 ;
        RECT 276.450 72.485 276.620 72.655 ;
        RECT 144.685 71.920 144.855 72.090 ;
        RECT 144.685 71.560 144.855 71.730 ;
        RECT 144.685 71.200 144.855 71.370 ;
        RECT 144.685 70.840 144.855 71.010 ;
        RECT 144.685 70.480 144.855 70.650 ;
        RECT 144.685 70.120 144.855 70.290 ;
        RECT 144.685 69.760 144.855 69.930 ;
        RECT 144.685 69.400 144.855 69.570 ;
        RECT 144.685 69.040 144.855 69.210 ;
        RECT 144.685 68.680 144.855 68.850 ;
        RECT 144.685 68.320 144.855 68.490 ;
        RECT 144.685 67.960 144.855 68.130 ;
        RECT 144.685 67.600 144.855 67.770 ;
        RECT 144.685 67.240 144.855 67.410 ;
        RECT 144.685 66.880 144.855 67.050 ;
        RECT 198.260 71.905 198.430 72.075 ;
        RECT 198.260 71.545 198.430 71.715 ;
        RECT 198.260 71.185 198.430 71.355 ;
        RECT 198.260 70.825 198.430 70.995 ;
        RECT 198.260 70.465 198.430 70.635 ;
        RECT 198.260 70.105 198.430 70.275 ;
        RECT 198.260 69.745 198.430 69.915 ;
        RECT 198.260 69.385 198.430 69.555 ;
        RECT 198.260 69.025 198.430 69.195 ;
        RECT 198.260 68.665 198.430 68.835 ;
        RECT 198.260 68.305 198.430 68.475 ;
        RECT 198.260 67.945 198.430 68.115 ;
        RECT 198.260 67.585 198.430 67.755 ;
        RECT 198.260 67.225 198.430 67.395 ;
        RECT 144.685 66.520 144.855 66.690 ;
        RECT 147.255 66.650 147.425 66.820 ;
        RECT 147.615 66.650 147.785 66.820 ;
        RECT 147.975 66.650 148.145 66.820 ;
        RECT 148.335 66.650 148.505 66.820 ;
        RECT 148.695 66.650 148.865 66.820 ;
        RECT 149.055 66.650 149.225 66.820 ;
        RECT 198.260 66.865 198.430 67.035 ;
        RECT 144.685 66.160 144.855 66.330 ;
        RECT 144.685 65.800 144.855 65.970 ;
        RECT 144.685 65.440 144.855 65.610 ;
        RECT 198.260 66.505 198.430 66.675 ;
        RECT 198.260 66.145 198.430 66.315 ;
        RECT 198.260 65.785 198.430 65.955 ;
        RECT 198.260 65.425 198.430 65.595 ;
        RECT 198.260 65.065 198.430 65.235 ;
        RECT 222.945 72.140 223.115 72.310 ;
        RECT 222.945 71.780 223.115 71.950 ;
        RECT 222.945 71.420 223.115 71.590 ;
        RECT 222.945 71.060 223.115 71.230 ;
        RECT 222.945 70.700 223.115 70.870 ;
        RECT 222.945 70.340 223.115 70.510 ;
        RECT 222.945 69.980 223.115 70.150 ;
        RECT 222.945 69.620 223.115 69.790 ;
        RECT 222.945 69.260 223.115 69.430 ;
        RECT 222.945 68.900 223.115 69.070 ;
        RECT 222.945 68.540 223.115 68.710 ;
        RECT 222.945 68.180 223.115 68.350 ;
        RECT 222.945 67.820 223.115 67.990 ;
        RECT 222.945 67.460 223.115 67.630 ;
        RECT 222.945 67.100 223.115 67.270 ;
        RECT 222.945 66.740 223.115 66.910 ;
        RECT 222.945 66.380 223.115 66.550 ;
        RECT 222.945 66.020 223.115 66.190 ;
        RECT 222.945 65.660 223.115 65.830 ;
        RECT 222.945 65.300 223.115 65.470 ;
        RECT 276.450 72.125 276.620 72.295 ;
        RECT 276.450 71.765 276.620 71.935 ;
        RECT 276.450 71.405 276.620 71.575 ;
        RECT 276.450 71.045 276.620 71.215 ;
        RECT 276.450 70.685 276.620 70.855 ;
        RECT 276.450 70.325 276.620 70.495 ;
        RECT 276.450 69.965 276.620 70.135 ;
        RECT 276.450 69.605 276.620 69.775 ;
        RECT 276.450 69.245 276.620 69.415 ;
        RECT 276.450 68.885 276.620 69.055 ;
        RECT 276.450 68.525 276.620 68.695 ;
        RECT 276.450 68.165 276.620 68.335 ;
        RECT 276.450 67.805 276.620 67.975 ;
        RECT 276.450 67.445 276.620 67.615 ;
        RECT 276.450 67.085 276.620 67.255 ;
        RECT 276.450 66.725 276.620 66.895 ;
        RECT 276.450 66.365 276.620 66.535 ;
        RECT 276.450 66.005 276.620 66.175 ;
        RECT 276.450 65.645 276.620 65.815 ;
        RECT 276.450 65.285 276.620 65.455 ;
        RECT 147.250 64.370 147.420 64.540 ;
        RECT 147.610 64.370 147.780 64.540 ;
        RECT 147.970 64.370 148.140 64.540 ;
        RECT 148.330 64.370 148.500 64.540 ;
        RECT 148.690 64.370 148.860 64.540 ;
        RECT 149.050 64.370 149.220 64.540 ;
        RECT 151.285 64.355 151.455 64.525 ;
        RECT 151.645 64.355 151.815 64.525 ;
        RECT 152.005 64.355 152.175 64.525 ;
        RECT 152.365 64.355 152.535 64.525 ;
        RECT 152.725 64.355 152.895 64.525 ;
        RECT 153.085 64.355 153.255 64.525 ;
        RECT 153.445 64.355 153.615 64.525 ;
        RECT 153.805 64.355 153.975 64.525 ;
        RECT 154.165 64.355 154.335 64.525 ;
        RECT 154.525 64.355 154.695 64.525 ;
        RECT 154.885 64.355 155.055 64.525 ;
        RECT 155.245 64.355 155.415 64.525 ;
        RECT 155.605 64.355 155.775 64.525 ;
        RECT 155.965 64.355 156.135 64.525 ;
        RECT 156.325 64.355 156.495 64.525 ;
        RECT 156.685 64.355 156.855 64.525 ;
        RECT 157.045 64.355 157.215 64.525 ;
        RECT 157.405 64.355 157.575 64.525 ;
        RECT 157.765 64.355 157.935 64.525 ;
        RECT 158.125 64.355 158.295 64.525 ;
        RECT 158.485 64.355 158.655 64.525 ;
        RECT 158.845 64.355 159.015 64.525 ;
        RECT 159.205 64.355 159.375 64.525 ;
        RECT 159.565 64.355 159.735 64.525 ;
        RECT 159.925 64.355 160.095 64.525 ;
        RECT 160.285 64.355 160.455 64.525 ;
        RECT 160.645 64.355 160.815 64.525 ;
        RECT 161.005 64.355 161.175 64.525 ;
        RECT 161.365 64.355 161.535 64.525 ;
        RECT 161.725 64.355 161.895 64.525 ;
        RECT 162.085 64.355 162.255 64.525 ;
        RECT 162.445 64.355 162.615 64.525 ;
        RECT 162.805 64.355 162.975 64.525 ;
        RECT 163.165 64.355 163.335 64.525 ;
        RECT 163.525 64.355 163.695 64.525 ;
        RECT 163.885 64.355 164.055 64.525 ;
        RECT 164.245 64.355 164.415 64.525 ;
        RECT 164.605 64.355 164.775 64.525 ;
        RECT 164.965 64.355 165.135 64.525 ;
        RECT 165.325 64.355 165.495 64.525 ;
        RECT 165.685 64.355 165.855 64.525 ;
        RECT 166.045 64.355 166.215 64.525 ;
        RECT 166.405 64.355 166.575 64.525 ;
        RECT 166.765 64.355 166.935 64.525 ;
        RECT 167.125 64.355 167.295 64.525 ;
        RECT 167.485 64.355 167.655 64.525 ;
        RECT 167.845 64.355 168.015 64.525 ;
        RECT 168.205 64.355 168.375 64.525 ;
        RECT 168.565 64.355 168.735 64.525 ;
        RECT 168.925 64.355 169.095 64.525 ;
        RECT 169.285 64.355 169.455 64.525 ;
        RECT 169.645 64.355 169.815 64.525 ;
        RECT 170.005 64.355 170.175 64.525 ;
        RECT 170.365 64.355 170.535 64.525 ;
        RECT 170.725 64.355 170.895 64.525 ;
        RECT 172.755 64.365 172.925 64.535 ;
        RECT 173.115 64.365 173.285 64.535 ;
        RECT 173.475 64.365 173.645 64.535 ;
        RECT 173.835 64.365 174.005 64.535 ;
        RECT 174.195 64.365 174.365 64.535 ;
        RECT 174.555 64.365 174.725 64.535 ;
        RECT 174.915 64.365 175.085 64.535 ;
        RECT 175.275 64.365 175.445 64.535 ;
        RECT 175.635 64.365 175.805 64.535 ;
        RECT 175.995 64.365 176.165 64.535 ;
        RECT 176.355 64.365 176.525 64.535 ;
        RECT 176.715 64.365 176.885 64.535 ;
        RECT 177.075 64.365 177.245 64.535 ;
        RECT 177.435 64.365 177.605 64.535 ;
        RECT 177.795 64.365 177.965 64.535 ;
        RECT 178.155 64.365 178.325 64.535 ;
        RECT 178.515 64.365 178.685 64.535 ;
        RECT 178.875 64.365 179.045 64.535 ;
        RECT 179.235 64.365 179.405 64.535 ;
        RECT 179.595 64.365 179.765 64.535 ;
        RECT 179.955 64.365 180.125 64.535 ;
        RECT 180.315 64.365 180.485 64.535 ;
        RECT 180.675 64.365 180.845 64.535 ;
        RECT 181.035 64.365 181.205 64.535 ;
        RECT 181.395 64.365 181.565 64.535 ;
        RECT 181.755 64.365 181.925 64.535 ;
        RECT 182.115 64.365 182.285 64.535 ;
        RECT 182.475 64.365 182.645 64.535 ;
        RECT 182.835 64.365 183.005 64.535 ;
        RECT 183.195 64.365 183.365 64.535 ;
        RECT 183.555 64.365 183.725 64.535 ;
        RECT 183.915 64.365 184.085 64.535 ;
        RECT 184.275 64.365 184.445 64.535 ;
        RECT 184.635 64.365 184.805 64.535 ;
        RECT 184.995 64.365 185.165 64.535 ;
        RECT 185.355 64.365 185.525 64.535 ;
        RECT 185.715 64.365 185.885 64.535 ;
        RECT 186.075 64.365 186.245 64.535 ;
        RECT 186.435 64.365 186.605 64.535 ;
        RECT 186.795 64.365 186.965 64.535 ;
        RECT 187.155 64.365 187.325 64.535 ;
        RECT 187.515 64.365 187.685 64.535 ;
        RECT 187.875 64.365 188.045 64.535 ;
        RECT 188.235 64.365 188.405 64.535 ;
        RECT 188.595 64.365 188.765 64.535 ;
        RECT 188.955 64.365 189.125 64.535 ;
        RECT 189.315 64.365 189.485 64.535 ;
        RECT 189.675 64.365 189.845 64.535 ;
        RECT 190.035 64.365 190.205 64.535 ;
        RECT 190.395 64.365 190.565 64.535 ;
        RECT 190.755 64.365 190.925 64.535 ;
        RECT 191.115 64.365 191.285 64.535 ;
        RECT 191.475 64.365 191.645 64.535 ;
        RECT 191.835 64.365 192.005 64.535 ;
        RECT 192.195 64.365 192.365 64.535 ;
        RECT 193.310 64.375 193.480 64.545 ;
        RECT 193.670 64.375 193.840 64.545 ;
        RECT 194.030 64.375 194.200 64.545 ;
        RECT 194.390 64.375 194.560 64.545 ;
        RECT 194.750 64.375 194.920 64.545 ;
        RECT 195.110 64.375 195.280 64.545 ;
        RECT 195.470 64.375 195.640 64.545 ;
        RECT 195.830 64.375 196.000 64.545 ;
        RECT 196.190 64.375 196.360 64.545 ;
        RECT 196.550 64.375 196.720 64.545 ;
        RECT 196.910 64.375 197.080 64.545 ;
        RECT 197.270 64.375 197.440 64.545 ;
        RECT 197.630 64.375 197.800 64.545 ;
        RECT 276.450 64.925 276.620 65.095 ;
        RECT 223.875 64.425 224.045 64.595 ;
        RECT 224.235 64.425 224.405 64.595 ;
        RECT 224.595 64.425 224.765 64.595 ;
        RECT 224.955 64.425 225.125 64.595 ;
        RECT 225.315 64.425 225.485 64.595 ;
        RECT 225.675 64.425 225.845 64.595 ;
        RECT 226.035 64.425 226.205 64.595 ;
        RECT 226.395 64.425 226.565 64.595 ;
        RECT 226.755 64.425 226.925 64.595 ;
        RECT 227.115 64.425 227.285 64.595 ;
        RECT 227.475 64.425 227.645 64.595 ;
        RECT 227.835 64.425 228.005 64.595 ;
        RECT 228.195 64.425 228.365 64.595 ;
        RECT 228.555 64.425 228.725 64.595 ;
        RECT 228.915 64.425 229.085 64.595 ;
        RECT 229.275 64.425 229.445 64.595 ;
        RECT 229.635 64.425 229.805 64.595 ;
        RECT 229.995 64.425 230.165 64.595 ;
        RECT 230.355 64.425 230.525 64.595 ;
        RECT 230.715 64.425 230.885 64.595 ;
        RECT 231.075 64.425 231.245 64.595 ;
        RECT 231.435 64.425 231.605 64.595 ;
        RECT 231.795 64.425 231.965 64.595 ;
        RECT 232.155 64.425 232.325 64.595 ;
        RECT 232.515 64.425 232.685 64.595 ;
        RECT 232.875 64.425 233.045 64.595 ;
        RECT 233.235 64.425 233.405 64.595 ;
        RECT 233.595 64.425 233.765 64.595 ;
        RECT 233.955 64.425 234.125 64.595 ;
        RECT 234.315 64.425 234.485 64.595 ;
        RECT 234.675 64.425 234.845 64.595 ;
        RECT 235.035 64.425 235.205 64.595 ;
        RECT 235.395 64.425 235.565 64.595 ;
        RECT 235.755 64.425 235.925 64.595 ;
        RECT 236.115 64.425 236.285 64.595 ;
        RECT 236.475 64.425 236.645 64.595 ;
        RECT 236.835 64.425 237.005 64.595 ;
        RECT 237.195 64.425 237.365 64.595 ;
        RECT 237.555 64.425 237.725 64.595 ;
        RECT 237.915 64.425 238.085 64.595 ;
        RECT 238.275 64.425 238.445 64.595 ;
        RECT 238.635 64.425 238.805 64.595 ;
        RECT 238.995 64.425 239.165 64.595 ;
        RECT 239.355 64.425 239.525 64.595 ;
        RECT 239.715 64.425 239.885 64.595 ;
        RECT 240.075 64.425 240.245 64.595 ;
        RECT 240.435 64.425 240.605 64.595 ;
        RECT 240.795 64.425 240.965 64.595 ;
        RECT 241.155 64.425 241.325 64.595 ;
        RECT 241.515 64.425 241.685 64.595 ;
        RECT 241.875 64.425 242.045 64.595 ;
        RECT 242.235 64.425 242.405 64.595 ;
        RECT 242.595 64.425 242.765 64.595 ;
        RECT 242.955 64.425 243.125 64.595 ;
        RECT 243.315 64.425 243.485 64.595 ;
        RECT 243.675 64.425 243.845 64.595 ;
        RECT 244.035 64.425 244.205 64.595 ;
        RECT 244.395 64.425 244.565 64.595 ;
        RECT 244.755 64.425 244.925 64.595 ;
        RECT 245.115 64.425 245.285 64.595 ;
        RECT 245.475 64.425 245.645 64.595 ;
        RECT 245.835 64.425 246.005 64.595 ;
        RECT 246.195 64.425 246.365 64.595 ;
        RECT 246.555 64.425 246.725 64.595 ;
        RECT 246.915 64.425 247.085 64.595 ;
        RECT 247.275 64.425 247.445 64.595 ;
        RECT 247.635 64.425 247.805 64.595 ;
        RECT 247.995 64.425 248.165 64.595 ;
        RECT 250.035 64.365 250.205 64.535 ;
        RECT 250.395 64.365 250.565 64.535 ;
        RECT 250.755 64.365 250.925 64.535 ;
        RECT 251.115 64.365 251.285 64.535 ;
        RECT 251.475 64.365 251.645 64.535 ;
        RECT 251.835 64.365 252.005 64.535 ;
        RECT 252.195 64.365 252.365 64.535 ;
        RECT 252.555 64.365 252.725 64.535 ;
        RECT 252.915 64.365 253.085 64.535 ;
        RECT 253.275 64.365 253.445 64.535 ;
        RECT 253.635 64.365 253.805 64.535 ;
        RECT 253.995 64.365 254.165 64.535 ;
        RECT 254.355 64.365 254.525 64.535 ;
        RECT 254.715 64.365 254.885 64.535 ;
        RECT 255.075 64.365 255.245 64.535 ;
        RECT 255.435 64.365 255.605 64.535 ;
        RECT 255.795 64.365 255.965 64.535 ;
        RECT 256.155 64.365 256.325 64.535 ;
        RECT 256.515 64.365 256.685 64.535 ;
        RECT 256.875 64.365 257.045 64.535 ;
        RECT 257.235 64.365 257.405 64.535 ;
        RECT 257.595 64.365 257.765 64.535 ;
        RECT 257.955 64.365 258.125 64.535 ;
        RECT 258.315 64.365 258.485 64.535 ;
        RECT 258.675 64.365 258.845 64.535 ;
        RECT 259.035 64.365 259.205 64.535 ;
        RECT 259.395 64.365 259.565 64.535 ;
        RECT 259.755 64.365 259.925 64.535 ;
        RECT 260.115 64.365 260.285 64.535 ;
        RECT 260.475 64.365 260.645 64.535 ;
        RECT 260.835 64.365 261.005 64.535 ;
        RECT 261.195 64.365 261.365 64.535 ;
        RECT 261.555 64.365 261.725 64.535 ;
        RECT 261.915 64.365 262.085 64.535 ;
        RECT 262.275 64.365 262.445 64.535 ;
        RECT 262.635 64.365 262.805 64.535 ;
        RECT 262.995 64.365 263.165 64.535 ;
        RECT 263.355 64.365 263.525 64.535 ;
        RECT 263.715 64.365 263.885 64.535 ;
        RECT 264.075 64.365 264.245 64.535 ;
        RECT 264.435 64.365 264.605 64.535 ;
        RECT 264.795 64.365 264.965 64.535 ;
        RECT 265.155 64.365 265.325 64.535 ;
        RECT 265.515 64.365 265.685 64.535 ;
        RECT 265.875 64.365 266.045 64.535 ;
        RECT 266.235 64.365 266.405 64.535 ;
        RECT 266.595 64.365 266.765 64.535 ;
        RECT 266.955 64.365 267.125 64.535 ;
        RECT 267.315 64.365 267.485 64.535 ;
        RECT 267.675 64.365 267.845 64.535 ;
        RECT 268.035 64.365 268.205 64.535 ;
        RECT 268.395 64.365 268.565 64.535 ;
        RECT 268.755 64.365 268.925 64.535 ;
        RECT 269.115 64.365 269.285 64.535 ;
        RECT 269.475 64.365 269.645 64.535 ;
      LAYER met1 ;
        RECT 151.000 133.210 220.010 134.030 ;
        RECT 249.865 133.800 269.770 133.815 ;
        RECT 249.865 133.795 274.205 133.800 ;
        RECT 249.805 133.365 274.205 133.795 ;
        RECT 249.805 133.360 269.830 133.365 ;
        RECT 249.865 133.340 269.770 133.360 ;
        RECT 144.350 65.070 145.085 131.540 ;
        RECT 271.995 131.200 274.155 133.365 ;
        RECT 206.045 96.635 206.510 99.285 ;
        RECT 205.990 96.065 207.170 96.245 ;
        RECT 205.990 95.955 207.265 96.065 ;
        RECT 204.925 95.725 207.265 95.955 ;
        RECT 204.925 95.590 205.345 95.725 ;
        RECT 205.990 95.630 207.265 95.725 ;
        RECT 205.990 95.330 207.170 95.630 ;
        RECT 206.015 92.860 207.195 93.090 ;
        RECT 206.005 92.750 207.260 92.860 ;
        RECT 204.930 92.740 207.260 92.750 ;
        RECT 204.925 92.520 207.260 92.740 ;
        RECT 204.925 92.510 205.345 92.520 ;
        RECT 206.005 92.425 207.260 92.520 ;
        RECT 206.015 92.175 207.195 92.425 ;
        RECT 206.055 89.855 207.235 90.075 ;
        RECT 206.010 89.765 207.265 89.855 ;
        RECT 204.940 89.660 207.265 89.765 ;
        RECT 204.925 89.535 207.265 89.660 ;
        RECT 204.925 89.430 205.345 89.535 ;
        RECT 206.010 89.420 207.265 89.535 ;
        RECT 206.055 89.160 207.235 89.420 ;
        RECT 200.235 84.230 200.705 85.820 ;
        RECT 204.925 85.605 205.345 85.790 ;
        RECT 206.045 85.715 207.225 85.955 ;
        RECT 206.020 85.605 207.275 85.715 ;
        RECT 207.955 85.605 208.375 85.790 ;
        RECT 204.925 85.560 208.410 85.605 ;
        RECT 204.945 85.360 208.410 85.560 ;
        RECT 206.020 85.280 207.275 85.360 ;
        RECT 206.045 85.040 207.225 85.280 ;
        RECT 208.910 79.740 212.670 80.370 ;
        RECT 208.325 78.480 208.745 78.510 ;
        RECT 208.320 78.220 208.750 78.480 ;
        RECT 209.655 78.220 211.925 79.740 ;
        RECT 212.835 78.480 213.255 78.510 ;
        RECT 212.830 78.220 213.260 78.480 ;
        RECT 208.320 76.330 213.260 78.220 ;
        RECT 208.320 76.010 208.750 76.330 ;
        RECT 208.325 75.990 208.745 76.010 ;
        RECT 209.655 74.740 211.925 76.330 ;
        RECT 212.830 76.010 213.260 76.330 ;
        RECT 212.835 75.990 213.255 76.010 ;
        RECT 209.060 74.110 212.520 74.740 ;
        RECT 209.135 73.520 212.515 74.110 ;
        RECT 197.605 73.515 223.215 73.520 ;
        RECT 197.605 72.395 223.265 73.515 ;
        RECT 147.155 65.070 149.315 66.910 ;
        RECT 197.605 65.070 198.710 72.395 ;
        RECT 144.345 63.965 198.710 65.070 ;
        RECT 222.510 64.835 223.265 72.395 ;
        RECT 275.970 64.835 276.985 133.975 ;
        RECT 222.510 64.080 276.985 64.835 ;
      LAYER via ;
        RECT 172.645 133.455 172.905 133.715 ;
        RECT 172.965 133.455 173.225 133.715 ;
        RECT 173.285 133.455 173.545 133.715 ;
        RECT 173.605 133.455 173.865 133.715 ;
        RECT 173.925 133.455 174.185 133.715 ;
        RECT 174.245 133.455 174.505 133.715 ;
        RECT 174.565 133.455 174.825 133.715 ;
        RECT 174.885 133.455 175.145 133.715 ;
        RECT 175.205 133.455 175.465 133.715 ;
        RECT 175.525 133.455 175.785 133.715 ;
        RECT 175.845 133.455 176.105 133.715 ;
        RECT 176.165 133.455 176.425 133.715 ;
        RECT 176.485 133.455 176.745 133.715 ;
        RECT 176.805 133.455 177.065 133.715 ;
        RECT 177.125 133.455 177.385 133.715 ;
        RECT 177.445 133.455 177.705 133.715 ;
        RECT 177.765 133.455 178.025 133.715 ;
        RECT 178.085 133.455 178.345 133.715 ;
        RECT 178.405 133.455 178.665 133.715 ;
        RECT 178.725 133.455 178.985 133.715 ;
        RECT 179.045 133.455 179.305 133.715 ;
        RECT 179.365 133.455 179.625 133.715 ;
        RECT 179.685 133.455 179.945 133.715 ;
        RECT 180.005 133.455 180.265 133.715 ;
        RECT 180.325 133.455 180.585 133.715 ;
        RECT 180.645 133.455 180.905 133.715 ;
        RECT 180.965 133.455 181.225 133.715 ;
        RECT 181.285 133.455 181.545 133.715 ;
        RECT 181.605 133.455 181.865 133.715 ;
        RECT 181.925 133.455 182.185 133.715 ;
        RECT 182.245 133.455 182.505 133.715 ;
        RECT 182.565 133.455 182.825 133.715 ;
        RECT 182.885 133.455 183.145 133.715 ;
        RECT 183.205 133.455 183.465 133.715 ;
        RECT 183.525 133.455 183.785 133.715 ;
        RECT 183.845 133.455 184.105 133.715 ;
        RECT 184.165 133.455 184.425 133.715 ;
        RECT 184.485 133.455 184.745 133.715 ;
        RECT 184.805 133.455 185.065 133.715 ;
        RECT 185.125 133.455 185.385 133.715 ;
        RECT 185.445 133.455 185.705 133.715 ;
        RECT 185.765 133.455 186.025 133.715 ;
        RECT 186.085 133.455 186.345 133.715 ;
        RECT 186.405 133.455 186.665 133.715 ;
        RECT 186.725 133.455 186.985 133.715 ;
        RECT 187.045 133.455 187.305 133.715 ;
        RECT 187.365 133.455 187.625 133.715 ;
        RECT 187.685 133.455 187.945 133.715 ;
        RECT 188.005 133.455 188.265 133.715 ;
        RECT 188.325 133.455 188.585 133.715 ;
        RECT 188.645 133.455 188.905 133.715 ;
        RECT 188.965 133.455 189.225 133.715 ;
        RECT 189.285 133.455 189.545 133.715 ;
        RECT 189.605 133.455 189.865 133.715 ;
        RECT 189.925 133.455 190.185 133.715 ;
        RECT 190.245 133.455 190.505 133.715 ;
        RECT 190.565 133.455 190.825 133.715 ;
        RECT 190.885 133.455 191.145 133.715 ;
        RECT 191.205 133.455 191.465 133.715 ;
        RECT 191.525 133.455 191.785 133.715 ;
        RECT 191.845 133.455 192.105 133.715 ;
        RECT 192.165 133.455 192.425 133.715 ;
        RECT 249.930 133.450 250.190 133.710 ;
        RECT 250.250 133.450 250.510 133.710 ;
        RECT 250.570 133.450 250.830 133.710 ;
        RECT 250.890 133.450 251.150 133.710 ;
        RECT 251.210 133.450 251.470 133.710 ;
        RECT 251.530 133.450 251.790 133.710 ;
        RECT 251.850 133.450 252.110 133.710 ;
        RECT 252.170 133.450 252.430 133.710 ;
        RECT 252.490 133.450 252.750 133.710 ;
        RECT 252.810 133.450 253.070 133.710 ;
        RECT 253.130 133.450 253.390 133.710 ;
        RECT 253.450 133.450 253.710 133.710 ;
        RECT 253.770 133.450 254.030 133.710 ;
        RECT 254.090 133.450 254.350 133.710 ;
        RECT 254.410 133.450 254.670 133.710 ;
        RECT 254.730 133.450 254.990 133.710 ;
        RECT 255.050 133.450 255.310 133.710 ;
        RECT 255.370 133.450 255.630 133.710 ;
        RECT 255.690 133.450 255.950 133.710 ;
        RECT 256.010 133.450 256.270 133.710 ;
        RECT 256.330 133.450 256.590 133.710 ;
        RECT 256.650 133.450 256.910 133.710 ;
        RECT 256.970 133.450 257.230 133.710 ;
        RECT 257.290 133.450 257.550 133.710 ;
        RECT 257.610 133.450 257.870 133.710 ;
        RECT 257.930 133.450 258.190 133.710 ;
        RECT 258.250 133.450 258.510 133.710 ;
        RECT 258.570 133.450 258.830 133.710 ;
        RECT 258.890 133.450 259.150 133.710 ;
        RECT 259.210 133.450 259.470 133.710 ;
        RECT 259.530 133.450 259.790 133.710 ;
        RECT 259.850 133.450 260.110 133.710 ;
        RECT 260.170 133.450 260.430 133.710 ;
        RECT 260.490 133.450 260.750 133.710 ;
        RECT 260.810 133.450 261.070 133.710 ;
        RECT 261.130 133.450 261.390 133.710 ;
        RECT 261.450 133.450 261.710 133.710 ;
        RECT 261.770 133.450 262.030 133.710 ;
        RECT 262.090 133.450 262.350 133.710 ;
        RECT 262.410 133.450 262.670 133.710 ;
        RECT 262.730 133.450 262.990 133.710 ;
        RECT 263.050 133.450 263.310 133.710 ;
        RECT 263.370 133.450 263.630 133.710 ;
        RECT 263.690 133.450 263.950 133.710 ;
        RECT 264.010 133.450 264.270 133.710 ;
        RECT 264.330 133.450 264.590 133.710 ;
        RECT 264.650 133.450 264.910 133.710 ;
        RECT 264.970 133.450 265.230 133.710 ;
        RECT 265.290 133.450 265.550 133.710 ;
        RECT 265.610 133.450 265.870 133.710 ;
        RECT 265.930 133.450 266.190 133.710 ;
        RECT 266.250 133.450 266.510 133.710 ;
        RECT 266.570 133.450 266.830 133.710 ;
        RECT 266.890 133.450 267.150 133.710 ;
        RECT 267.210 133.450 267.470 133.710 ;
        RECT 267.530 133.450 267.790 133.710 ;
        RECT 267.850 133.450 268.110 133.710 ;
        RECT 268.170 133.450 268.430 133.710 ;
        RECT 268.490 133.450 268.750 133.710 ;
        RECT 268.810 133.450 269.070 133.710 ;
        RECT 269.130 133.450 269.390 133.710 ;
        RECT 269.450 133.450 269.710 133.710 ;
        RECT 206.150 98.950 206.410 99.210 ;
        RECT 206.150 98.630 206.410 98.890 ;
        RECT 206.150 98.310 206.410 98.570 ;
        RECT 206.150 97.990 206.410 98.250 ;
        RECT 206.150 97.670 206.410 97.930 ;
        RECT 206.150 97.350 206.410 97.610 ;
        RECT 206.150 97.030 206.410 97.290 ;
        RECT 206.150 96.710 206.410 96.970 ;
        RECT 206.130 95.500 207.030 96.080 ;
        RECT 206.155 92.345 207.055 92.925 ;
        RECT 206.195 89.330 207.095 89.910 ;
        RECT 200.340 85.495 200.600 85.755 ;
        RECT 200.340 85.175 200.600 85.435 ;
        RECT 200.340 84.855 200.600 85.115 ;
        RECT 206.185 85.210 207.085 85.790 ;
        RECT 200.340 84.535 200.600 84.795 ;
        RECT 172.670 64.320 172.930 64.580 ;
        RECT 172.990 64.320 173.250 64.580 ;
        RECT 173.310 64.320 173.570 64.580 ;
        RECT 173.630 64.320 173.890 64.580 ;
        RECT 173.950 64.320 174.210 64.580 ;
        RECT 174.270 64.320 174.530 64.580 ;
        RECT 174.590 64.320 174.850 64.580 ;
        RECT 174.910 64.320 175.170 64.580 ;
        RECT 175.230 64.320 175.490 64.580 ;
        RECT 175.550 64.320 175.810 64.580 ;
        RECT 175.870 64.320 176.130 64.580 ;
        RECT 176.190 64.320 176.450 64.580 ;
        RECT 176.510 64.320 176.770 64.580 ;
        RECT 176.830 64.320 177.090 64.580 ;
        RECT 177.150 64.320 177.410 64.580 ;
        RECT 177.470 64.320 177.730 64.580 ;
        RECT 177.790 64.320 178.050 64.580 ;
        RECT 178.110 64.320 178.370 64.580 ;
        RECT 178.430 64.320 178.690 64.580 ;
        RECT 178.750 64.320 179.010 64.580 ;
        RECT 179.070 64.320 179.330 64.580 ;
        RECT 179.390 64.320 179.650 64.580 ;
        RECT 179.710 64.320 179.970 64.580 ;
        RECT 180.030 64.320 180.290 64.580 ;
        RECT 180.350 64.320 180.610 64.580 ;
        RECT 180.670 64.320 180.930 64.580 ;
        RECT 180.990 64.320 181.250 64.580 ;
        RECT 181.310 64.320 181.570 64.580 ;
        RECT 181.630 64.320 181.890 64.580 ;
        RECT 181.950 64.320 182.210 64.580 ;
        RECT 182.270 64.320 182.530 64.580 ;
        RECT 182.590 64.320 182.850 64.580 ;
        RECT 182.910 64.320 183.170 64.580 ;
        RECT 183.230 64.320 183.490 64.580 ;
        RECT 183.550 64.320 183.810 64.580 ;
        RECT 183.870 64.320 184.130 64.580 ;
        RECT 184.190 64.320 184.450 64.580 ;
        RECT 184.510 64.320 184.770 64.580 ;
        RECT 184.830 64.320 185.090 64.580 ;
        RECT 185.150 64.320 185.410 64.580 ;
        RECT 185.470 64.320 185.730 64.580 ;
        RECT 185.790 64.320 186.050 64.580 ;
        RECT 186.110 64.320 186.370 64.580 ;
        RECT 186.430 64.320 186.690 64.580 ;
        RECT 186.750 64.320 187.010 64.580 ;
        RECT 187.070 64.320 187.330 64.580 ;
        RECT 187.390 64.320 187.650 64.580 ;
        RECT 187.710 64.320 187.970 64.580 ;
        RECT 188.030 64.320 188.290 64.580 ;
        RECT 188.350 64.320 188.610 64.580 ;
        RECT 188.670 64.320 188.930 64.580 ;
        RECT 188.990 64.320 189.250 64.580 ;
        RECT 189.310 64.320 189.570 64.580 ;
        RECT 189.630 64.320 189.890 64.580 ;
        RECT 189.950 64.320 190.210 64.580 ;
        RECT 190.270 64.320 190.530 64.580 ;
        RECT 190.590 64.320 190.850 64.580 ;
        RECT 190.910 64.320 191.170 64.580 ;
        RECT 191.230 64.320 191.490 64.580 ;
        RECT 191.550 64.320 191.810 64.580 ;
        RECT 191.870 64.320 192.130 64.580 ;
        RECT 192.190 64.320 192.450 64.580 ;
        RECT 249.950 64.320 250.210 64.580 ;
        RECT 250.270 64.320 250.530 64.580 ;
        RECT 250.590 64.320 250.850 64.580 ;
        RECT 250.910 64.320 251.170 64.580 ;
        RECT 251.230 64.320 251.490 64.580 ;
        RECT 251.550 64.320 251.810 64.580 ;
        RECT 251.870 64.320 252.130 64.580 ;
        RECT 252.190 64.320 252.450 64.580 ;
        RECT 252.510 64.320 252.770 64.580 ;
        RECT 252.830 64.320 253.090 64.580 ;
        RECT 253.150 64.320 253.410 64.580 ;
        RECT 253.470 64.320 253.730 64.580 ;
        RECT 253.790 64.320 254.050 64.580 ;
        RECT 254.110 64.320 254.370 64.580 ;
        RECT 254.430 64.320 254.690 64.580 ;
        RECT 254.750 64.320 255.010 64.580 ;
        RECT 255.070 64.320 255.330 64.580 ;
        RECT 255.390 64.320 255.650 64.580 ;
        RECT 255.710 64.320 255.970 64.580 ;
        RECT 256.030 64.320 256.290 64.580 ;
        RECT 256.350 64.320 256.610 64.580 ;
        RECT 256.670 64.320 256.930 64.580 ;
        RECT 256.990 64.320 257.250 64.580 ;
        RECT 257.310 64.320 257.570 64.580 ;
        RECT 257.630 64.320 257.890 64.580 ;
        RECT 257.950 64.320 258.210 64.580 ;
        RECT 258.270 64.320 258.530 64.580 ;
        RECT 258.590 64.320 258.850 64.580 ;
        RECT 258.910 64.320 259.170 64.580 ;
        RECT 259.230 64.320 259.490 64.580 ;
        RECT 259.550 64.320 259.810 64.580 ;
        RECT 259.870 64.320 260.130 64.580 ;
        RECT 260.190 64.320 260.450 64.580 ;
        RECT 260.510 64.320 260.770 64.580 ;
        RECT 260.830 64.320 261.090 64.580 ;
        RECT 261.150 64.320 261.410 64.580 ;
        RECT 261.470 64.320 261.730 64.580 ;
        RECT 261.790 64.320 262.050 64.580 ;
        RECT 262.110 64.320 262.370 64.580 ;
        RECT 262.430 64.320 262.690 64.580 ;
        RECT 262.750 64.320 263.010 64.580 ;
        RECT 263.070 64.320 263.330 64.580 ;
        RECT 263.390 64.320 263.650 64.580 ;
        RECT 263.710 64.320 263.970 64.580 ;
        RECT 264.030 64.320 264.290 64.580 ;
        RECT 264.350 64.320 264.610 64.580 ;
        RECT 264.670 64.320 264.930 64.580 ;
        RECT 264.990 64.320 265.250 64.580 ;
        RECT 265.310 64.320 265.570 64.580 ;
        RECT 265.630 64.320 265.890 64.580 ;
        RECT 265.950 64.320 266.210 64.580 ;
        RECT 266.270 64.320 266.530 64.580 ;
        RECT 266.590 64.320 266.850 64.580 ;
        RECT 266.910 64.320 267.170 64.580 ;
        RECT 267.230 64.320 267.490 64.580 ;
        RECT 267.550 64.320 267.810 64.580 ;
        RECT 267.870 64.320 268.130 64.580 ;
        RECT 268.190 64.320 268.450 64.580 ;
        RECT 268.510 64.320 268.770 64.580 ;
        RECT 268.830 64.320 269.090 64.580 ;
        RECT 269.150 64.320 269.410 64.580 ;
        RECT 269.470 64.320 269.730 64.580 ;
      LAYER met2 ;
        RECT 172.525 100.810 192.525 134.100 ;
        RECT 249.825 133.765 269.825 134.100 ;
        RECT 249.815 133.390 269.825 133.765 ;
        RECT 172.525 94.780 207.680 100.810 ;
        RECT 172.525 89.925 192.525 94.780 ;
        RECT 205.445 89.925 207.680 94.780 ;
        RECT 172.525 84.530 207.680 89.925 ;
        RECT 172.525 83.895 198.490 84.530 ;
        RECT 172.525 63.930 192.525 83.895 ;
        RECT 249.825 63.930 269.825 133.390 ;
      LAYER via2 ;
        RECT 176.990 133.720 177.270 134.000 ;
        RECT 177.390 133.720 177.670 134.000 ;
        RECT 177.790 133.720 178.070 134.000 ;
        RECT 178.190 133.720 178.470 134.000 ;
        RECT 180.320 133.720 180.600 134.000 ;
        RECT 180.720 133.720 181.000 134.000 ;
        RECT 181.120 133.720 181.400 134.000 ;
        RECT 181.520 133.720 181.800 134.000 ;
        RECT 183.615 133.700 183.895 133.980 ;
        RECT 184.015 133.700 184.295 133.980 ;
        RECT 184.415 133.700 184.695 133.980 ;
        RECT 184.815 133.700 185.095 133.980 ;
        RECT 186.930 133.700 187.210 133.980 ;
        RECT 187.330 133.700 187.610 133.980 ;
        RECT 187.730 133.700 188.010 133.980 ;
        RECT 188.130 133.700 188.410 133.980 ;
        RECT 176.990 133.160 177.270 133.440 ;
        RECT 177.390 133.160 177.670 133.440 ;
        RECT 177.790 133.160 178.070 133.440 ;
        RECT 178.190 133.160 178.470 133.440 ;
        RECT 180.320 133.160 180.600 133.440 ;
        RECT 180.720 133.160 181.000 133.440 ;
        RECT 181.120 133.160 181.400 133.440 ;
        RECT 181.520 133.160 181.800 133.440 ;
        RECT 183.615 133.140 183.895 133.420 ;
        RECT 184.015 133.140 184.295 133.420 ;
        RECT 184.415 133.140 184.695 133.420 ;
        RECT 184.815 133.140 185.095 133.420 ;
        RECT 186.930 133.140 187.210 133.420 ;
        RECT 187.330 133.140 187.610 133.420 ;
        RECT 187.730 133.140 188.010 133.420 ;
        RECT 188.130 133.140 188.410 133.420 ;
        RECT 254.175 133.720 254.455 134.000 ;
        RECT 254.575 133.720 254.855 134.000 ;
        RECT 254.975 133.720 255.255 134.000 ;
        RECT 255.375 133.720 255.655 134.000 ;
        RECT 257.505 133.720 257.785 134.000 ;
        RECT 257.905 133.720 258.185 134.000 ;
        RECT 258.305 133.720 258.585 134.000 ;
        RECT 258.705 133.720 258.985 134.000 ;
        RECT 260.800 133.700 261.080 133.980 ;
        RECT 261.200 133.700 261.480 133.980 ;
        RECT 261.600 133.700 261.880 133.980 ;
        RECT 262.000 133.700 262.280 133.980 ;
        RECT 264.115 133.700 264.395 133.980 ;
        RECT 264.515 133.700 264.795 133.980 ;
        RECT 264.915 133.700 265.195 133.980 ;
        RECT 265.315 133.700 265.595 133.980 ;
        RECT 176.990 132.565 177.270 132.845 ;
        RECT 177.390 132.565 177.670 132.845 ;
        RECT 177.790 132.565 178.070 132.845 ;
        RECT 178.190 132.565 178.470 132.845 ;
        RECT 180.320 132.565 180.600 132.845 ;
        RECT 180.720 132.565 181.000 132.845 ;
        RECT 181.120 132.565 181.400 132.845 ;
        RECT 181.520 132.565 181.800 132.845 ;
        RECT 183.615 132.545 183.895 132.825 ;
        RECT 184.015 132.545 184.295 132.825 ;
        RECT 184.415 132.545 184.695 132.825 ;
        RECT 184.815 132.545 185.095 132.825 ;
        RECT 186.930 132.545 187.210 132.825 ;
        RECT 187.330 132.545 187.610 132.825 ;
        RECT 187.730 132.545 188.010 132.825 ;
        RECT 188.130 132.545 188.410 132.825 ;
        RECT 254.175 133.160 254.455 133.440 ;
        RECT 254.575 133.160 254.855 133.440 ;
        RECT 254.975 133.160 255.255 133.440 ;
        RECT 255.375 133.160 255.655 133.440 ;
        RECT 257.505 133.160 257.785 133.440 ;
        RECT 257.905 133.160 258.185 133.440 ;
        RECT 258.305 133.160 258.585 133.440 ;
        RECT 258.705 133.160 258.985 133.440 ;
        RECT 260.800 133.140 261.080 133.420 ;
        RECT 261.200 133.140 261.480 133.420 ;
        RECT 261.600 133.140 261.880 133.420 ;
        RECT 262.000 133.140 262.280 133.420 ;
        RECT 264.115 133.140 264.395 133.420 ;
        RECT 264.515 133.140 264.795 133.420 ;
        RECT 264.915 133.140 265.195 133.420 ;
        RECT 265.315 133.140 265.595 133.420 ;
        RECT 254.175 132.565 254.455 132.845 ;
        RECT 254.575 132.565 254.855 132.845 ;
        RECT 254.975 132.565 255.255 132.845 ;
        RECT 255.375 132.565 255.655 132.845 ;
        RECT 257.505 132.565 257.785 132.845 ;
        RECT 257.905 132.565 258.185 132.845 ;
        RECT 258.305 132.565 258.585 132.845 ;
        RECT 258.705 132.565 258.985 132.845 ;
        RECT 260.800 132.545 261.080 132.825 ;
        RECT 261.200 132.545 261.480 132.825 ;
        RECT 261.600 132.545 261.880 132.825 ;
        RECT 262.000 132.545 262.280 132.825 ;
        RECT 264.115 132.545 264.395 132.825 ;
        RECT 264.515 132.545 264.795 132.825 ;
        RECT 264.915 132.545 265.195 132.825 ;
        RECT 265.315 132.545 265.595 132.825 ;
        RECT 176.990 65.260 177.270 65.540 ;
        RECT 177.390 65.260 177.670 65.540 ;
        RECT 177.790 65.260 178.070 65.540 ;
        RECT 178.190 65.260 178.470 65.540 ;
        RECT 180.320 65.260 180.600 65.540 ;
        RECT 180.720 65.260 181.000 65.540 ;
        RECT 181.120 65.260 181.400 65.540 ;
        RECT 181.520 65.260 181.800 65.540 ;
        RECT 183.615 65.240 183.895 65.520 ;
        RECT 184.015 65.240 184.295 65.520 ;
        RECT 184.415 65.240 184.695 65.520 ;
        RECT 184.815 65.240 185.095 65.520 ;
        RECT 186.930 65.240 187.210 65.520 ;
        RECT 187.330 65.240 187.610 65.520 ;
        RECT 187.730 65.240 188.010 65.520 ;
        RECT 188.130 65.240 188.410 65.520 ;
        RECT 176.990 64.700 177.270 64.980 ;
        RECT 177.390 64.700 177.670 64.980 ;
        RECT 177.790 64.700 178.070 64.980 ;
        RECT 178.190 64.700 178.470 64.980 ;
        RECT 180.320 64.700 180.600 64.980 ;
        RECT 180.720 64.700 181.000 64.980 ;
        RECT 181.120 64.700 181.400 64.980 ;
        RECT 181.520 64.700 181.800 64.980 ;
        RECT 183.615 64.680 183.895 64.960 ;
        RECT 184.015 64.680 184.295 64.960 ;
        RECT 184.415 64.680 184.695 64.960 ;
        RECT 184.815 64.680 185.095 64.960 ;
        RECT 186.930 64.680 187.210 64.960 ;
        RECT 187.330 64.680 187.610 64.960 ;
        RECT 187.730 64.680 188.010 64.960 ;
        RECT 188.130 64.680 188.410 64.960 ;
        RECT 176.990 64.105 177.270 64.385 ;
        RECT 177.390 64.105 177.670 64.385 ;
        RECT 177.790 64.105 178.070 64.385 ;
        RECT 178.190 64.105 178.470 64.385 ;
        RECT 180.320 64.105 180.600 64.385 ;
        RECT 180.720 64.105 181.000 64.385 ;
        RECT 181.120 64.105 181.400 64.385 ;
        RECT 181.520 64.105 181.800 64.385 ;
        RECT 183.615 64.085 183.895 64.365 ;
        RECT 184.015 64.085 184.295 64.365 ;
        RECT 184.415 64.085 184.695 64.365 ;
        RECT 184.815 64.085 185.095 64.365 ;
        RECT 186.930 64.085 187.210 64.365 ;
        RECT 187.330 64.085 187.610 64.365 ;
        RECT 187.730 64.085 188.010 64.365 ;
        RECT 188.130 64.085 188.410 64.365 ;
        RECT 254.175 65.260 254.455 65.540 ;
        RECT 254.575 65.260 254.855 65.540 ;
        RECT 254.975 65.260 255.255 65.540 ;
        RECT 255.375 65.260 255.655 65.540 ;
        RECT 257.505 65.260 257.785 65.540 ;
        RECT 257.905 65.260 258.185 65.540 ;
        RECT 258.305 65.260 258.585 65.540 ;
        RECT 258.705 65.260 258.985 65.540 ;
        RECT 260.800 65.240 261.080 65.520 ;
        RECT 261.200 65.240 261.480 65.520 ;
        RECT 261.600 65.240 261.880 65.520 ;
        RECT 262.000 65.240 262.280 65.520 ;
        RECT 264.115 65.240 264.395 65.520 ;
        RECT 264.515 65.240 264.795 65.520 ;
        RECT 264.915 65.240 265.195 65.520 ;
        RECT 265.315 65.240 265.595 65.520 ;
        RECT 254.175 64.700 254.455 64.980 ;
        RECT 254.575 64.700 254.855 64.980 ;
        RECT 254.975 64.700 255.255 64.980 ;
        RECT 255.375 64.700 255.655 64.980 ;
        RECT 257.505 64.700 257.785 64.980 ;
        RECT 257.905 64.700 258.185 64.980 ;
        RECT 258.305 64.700 258.585 64.980 ;
        RECT 258.705 64.700 258.985 64.980 ;
        RECT 260.800 64.680 261.080 64.960 ;
        RECT 261.200 64.680 261.480 64.960 ;
        RECT 261.600 64.680 261.880 64.960 ;
        RECT 262.000 64.680 262.280 64.960 ;
        RECT 264.115 64.680 264.395 64.960 ;
        RECT 264.515 64.680 264.795 64.960 ;
        RECT 264.915 64.680 265.195 64.960 ;
        RECT 265.315 64.680 265.595 64.960 ;
        RECT 254.175 64.105 254.455 64.385 ;
        RECT 254.575 64.105 254.855 64.385 ;
        RECT 254.975 64.105 255.255 64.385 ;
        RECT 255.375 64.105 255.655 64.385 ;
        RECT 257.505 64.105 257.785 64.385 ;
        RECT 257.905 64.105 258.185 64.385 ;
        RECT 258.305 64.105 258.585 64.385 ;
        RECT 258.705 64.105 258.985 64.385 ;
        RECT 260.800 64.085 261.080 64.365 ;
        RECT 261.200 64.085 261.480 64.365 ;
        RECT 261.600 64.085 261.880 64.365 ;
        RECT 262.000 64.085 262.280 64.365 ;
        RECT 264.115 64.085 264.395 64.365 ;
        RECT 264.515 64.085 264.795 64.365 ;
        RECT 264.915 64.085 265.195 64.365 ;
        RECT 265.315 64.085 265.595 64.365 ;
      LAYER met3 ;
        RECT 172.525 132.390 192.525 134.100 ;
        RECT 249.710 132.390 269.710 134.100 ;
        RECT 172.525 63.930 192.525 65.640 ;
        RECT 249.710 63.930 269.710 65.640 ;
      LAYER via3 ;
        RECT 176.970 133.700 177.290 134.020 ;
        RECT 177.370 133.700 177.690 134.020 ;
        RECT 177.770 133.700 178.090 134.020 ;
        RECT 178.170 133.700 178.490 134.020 ;
        RECT 180.300 133.700 180.620 134.020 ;
        RECT 180.700 133.700 181.020 134.020 ;
        RECT 181.100 133.700 181.420 134.020 ;
        RECT 181.500 133.700 181.820 134.020 ;
        RECT 183.595 133.680 183.915 134.000 ;
        RECT 183.995 133.680 184.315 134.000 ;
        RECT 184.395 133.680 184.715 134.000 ;
        RECT 184.795 133.680 185.115 134.000 ;
        RECT 186.910 133.680 187.230 134.000 ;
        RECT 187.310 133.680 187.630 134.000 ;
        RECT 187.710 133.680 188.030 134.000 ;
        RECT 188.110 133.680 188.430 134.000 ;
        RECT 176.970 133.140 177.290 133.460 ;
        RECT 177.370 133.140 177.690 133.460 ;
        RECT 177.770 133.140 178.090 133.460 ;
        RECT 178.170 133.140 178.490 133.460 ;
        RECT 180.300 133.140 180.620 133.460 ;
        RECT 180.700 133.140 181.020 133.460 ;
        RECT 181.100 133.140 181.420 133.460 ;
        RECT 181.500 133.140 181.820 133.460 ;
        RECT 183.595 133.120 183.915 133.440 ;
        RECT 183.995 133.120 184.315 133.440 ;
        RECT 184.395 133.120 184.715 133.440 ;
        RECT 184.795 133.120 185.115 133.440 ;
        RECT 186.910 133.120 187.230 133.440 ;
        RECT 187.310 133.120 187.630 133.440 ;
        RECT 187.710 133.120 188.030 133.440 ;
        RECT 188.110 133.120 188.430 133.440 ;
        RECT 176.970 132.545 177.290 132.865 ;
        RECT 177.370 132.545 177.690 132.865 ;
        RECT 177.770 132.545 178.090 132.865 ;
        RECT 178.170 132.545 178.490 132.865 ;
        RECT 180.300 132.545 180.620 132.865 ;
        RECT 180.700 132.545 181.020 132.865 ;
        RECT 181.100 132.545 181.420 132.865 ;
        RECT 181.500 132.545 181.820 132.865 ;
        RECT 183.595 132.525 183.915 132.845 ;
        RECT 183.995 132.525 184.315 132.845 ;
        RECT 184.395 132.525 184.715 132.845 ;
        RECT 184.795 132.525 185.115 132.845 ;
        RECT 186.910 132.525 187.230 132.845 ;
        RECT 187.310 132.525 187.630 132.845 ;
        RECT 187.710 132.525 188.030 132.845 ;
        RECT 188.110 132.525 188.430 132.845 ;
        RECT 254.155 133.700 254.475 134.020 ;
        RECT 254.555 133.700 254.875 134.020 ;
        RECT 254.955 133.700 255.275 134.020 ;
        RECT 255.355 133.700 255.675 134.020 ;
        RECT 257.485 133.700 257.805 134.020 ;
        RECT 257.885 133.700 258.205 134.020 ;
        RECT 258.285 133.700 258.605 134.020 ;
        RECT 258.685 133.700 259.005 134.020 ;
        RECT 260.780 133.680 261.100 134.000 ;
        RECT 261.180 133.680 261.500 134.000 ;
        RECT 261.580 133.680 261.900 134.000 ;
        RECT 261.980 133.680 262.300 134.000 ;
        RECT 264.095 133.680 264.415 134.000 ;
        RECT 264.495 133.680 264.815 134.000 ;
        RECT 264.895 133.680 265.215 134.000 ;
        RECT 265.295 133.680 265.615 134.000 ;
        RECT 254.155 133.140 254.475 133.460 ;
        RECT 254.555 133.140 254.875 133.460 ;
        RECT 254.955 133.140 255.275 133.460 ;
        RECT 255.355 133.140 255.675 133.460 ;
        RECT 257.485 133.140 257.805 133.460 ;
        RECT 257.885 133.140 258.205 133.460 ;
        RECT 258.285 133.140 258.605 133.460 ;
        RECT 258.685 133.140 259.005 133.460 ;
        RECT 260.780 133.120 261.100 133.440 ;
        RECT 261.180 133.120 261.500 133.440 ;
        RECT 261.580 133.120 261.900 133.440 ;
        RECT 261.980 133.120 262.300 133.440 ;
        RECT 264.095 133.120 264.415 133.440 ;
        RECT 264.495 133.120 264.815 133.440 ;
        RECT 264.895 133.120 265.215 133.440 ;
        RECT 265.295 133.120 265.615 133.440 ;
        RECT 254.155 132.545 254.475 132.865 ;
        RECT 254.555 132.545 254.875 132.865 ;
        RECT 254.955 132.545 255.275 132.865 ;
        RECT 255.355 132.545 255.675 132.865 ;
        RECT 257.485 132.545 257.805 132.865 ;
        RECT 257.885 132.545 258.205 132.865 ;
        RECT 258.285 132.545 258.605 132.865 ;
        RECT 258.685 132.545 259.005 132.865 ;
        RECT 260.780 132.525 261.100 132.845 ;
        RECT 261.180 132.525 261.500 132.845 ;
        RECT 261.580 132.525 261.900 132.845 ;
        RECT 261.980 132.525 262.300 132.845 ;
        RECT 264.095 132.525 264.415 132.845 ;
        RECT 264.495 132.525 264.815 132.845 ;
        RECT 264.895 132.525 265.215 132.845 ;
        RECT 265.295 132.525 265.615 132.845 ;
        RECT 176.970 65.240 177.290 65.560 ;
        RECT 177.370 65.240 177.690 65.560 ;
        RECT 177.770 65.240 178.090 65.560 ;
        RECT 178.170 65.240 178.490 65.560 ;
        RECT 180.300 65.240 180.620 65.560 ;
        RECT 180.700 65.240 181.020 65.560 ;
        RECT 181.100 65.240 181.420 65.560 ;
        RECT 181.500 65.240 181.820 65.560 ;
        RECT 183.595 65.220 183.915 65.540 ;
        RECT 183.995 65.220 184.315 65.540 ;
        RECT 184.395 65.220 184.715 65.540 ;
        RECT 184.795 65.220 185.115 65.540 ;
        RECT 186.910 65.220 187.230 65.540 ;
        RECT 187.310 65.220 187.630 65.540 ;
        RECT 187.710 65.220 188.030 65.540 ;
        RECT 188.110 65.220 188.430 65.540 ;
        RECT 176.970 64.680 177.290 65.000 ;
        RECT 177.370 64.680 177.690 65.000 ;
        RECT 177.770 64.680 178.090 65.000 ;
        RECT 178.170 64.680 178.490 65.000 ;
        RECT 180.300 64.680 180.620 65.000 ;
        RECT 180.700 64.680 181.020 65.000 ;
        RECT 181.100 64.680 181.420 65.000 ;
        RECT 181.500 64.680 181.820 65.000 ;
        RECT 183.595 64.660 183.915 64.980 ;
        RECT 183.995 64.660 184.315 64.980 ;
        RECT 184.395 64.660 184.715 64.980 ;
        RECT 184.795 64.660 185.115 64.980 ;
        RECT 186.910 64.660 187.230 64.980 ;
        RECT 187.310 64.660 187.630 64.980 ;
        RECT 187.710 64.660 188.030 64.980 ;
        RECT 188.110 64.660 188.430 64.980 ;
        RECT 176.970 64.085 177.290 64.405 ;
        RECT 177.370 64.085 177.690 64.405 ;
        RECT 177.770 64.085 178.090 64.405 ;
        RECT 178.170 64.085 178.490 64.405 ;
        RECT 180.300 64.085 180.620 64.405 ;
        RECT 180.700 64.085 181.020 64.405 ;
        RECT 181.100 64.085 181.420 64.405 ;
        RECT 181.500 64.085 181.820 64.405 ;
        RECT 183.595 64.065 183.915 64.385 ;
        RECT 183.995 64.065 184.315 64.385 ;
        RECT 184.395 64.065 184.715 64.385 ;
        RECT 184.795 64.065 185.115 64.385 ;
        RECT 186.910 64.065 187.230 64.385 ;
        RECT 187.310 64.065 187.630 64.385 ;
        RECT 187.710 64.065 188.030 64.385 ;
        RECT 188.110 64.065 188.430 64.385 ;
        RECT 254.155 65.240 254.475 65.560 ;
        RECT 254.555 65.240 254.875 65.560 ;
        RECT 254.955 65.240 255.275 65.560 ;
        RECT 255.355 65.240 255.675 65.560 ;
        RECT 257.485 65.240 257.805 65.560 ;
        RECT 257.885 65.240 258.205 65.560 ;
        RECT 258.285 65.240 258.605 65.560 ;
        RECT 258.685 65.240 259.005 65.560 ;
        RECT 260.780 65.220 261.100 65.540 ;
        RECT 261.180 65.220 261.500 65.540 ;
        RECT 261.580 65.220 261.900 65.540 ;
        RECT 261.980 65.220 262.300 65.540 ;
        RECT 264.095 65.220 264.415 65.540 ;
        RECT 264.495 65.220 264.815 65.540 ;
        RECT 264.895 65.220 265.215 65.540 ;
        RECT 265.295 65.220 265.615 65.540 ;
        RECT 254.155 64.680 254.475 65.000 ;
        RECT 254.555 64.680 254.875 65.000 ;
        RECT 254.955 64.680 255.275 65.000 ;
        RECT 255.355 64.680 255.675 65.000 ;
        RECT 257.485 64.680 257.805 65.000 ;
        RECT 257.885 64.680 258.205 65.000 ;
        RECT 258.285 64.680 258.605 65.000 ;
        RECT 258.685 64.680 259.005 65.000 ;
        RECT 260.780 64.660 261.100 64.980 ;
        RECT 261.180 64.660 261.500 64.980 ;
        RECT 261.580 64.660 261.900 64.980 ;
        RECT 261.980 64.660 262.300 64.980 ;
        RECT 264.095 64.660 264.415 64.980 ;
        RECT 264.495 64.660 264.815 64.980 ;
        RECT 264.895 64.660 265.215 64.980 ;
        RECT 265.295 64.660 265.615 64.980 ;
        RECT 254.155 64.085 254.475 64.405 ;
        RECT 254.555 64.085 254.875 64.405 ;
        RECT 254.955 64.085 255.275 64.405 ;
        RECT 255.355 64.085 255.675 64.405 ;
        RECT 257.485 64.085 257.805 64.405 ;
        RECT 257.885 64.085 258.205 64.405 ;
        RECT 258.285 64.085 258.605 64.405 ;
        RECT 258.685 64.085 259.005 64.405 ;
        RECT 260.780 64.065 261.100 64.385 ;
        RECT 261.180 64.065 261.500 64.385 ;
        RECT 261.580 64.065 261.900 64.385 ;
        RECT 261.980 64.065 262.300 64.385 ;
        RECT 264.095 64.065 264.415 64.385 ;
        RECT 264.495 64.065 264.815 64.385 ;
        RECT 264.895 64.065 265.215 64.385 ;
        RECT 265.295 64.065 265.615 64.385 ;
      LAYER met4 ;
        RECT 176.935 3.300 178.535 211.800 ;
        RECT 180.235 3.300 181.835 211.800 ;
        RECT 183.535 3.300 185.135 211.800 ;
        RECT 186.835 3.300 188.435 211.800 ;
        RECT 254.120 3.300 255.720 211.800 ;
        RECT 257.420 3.300 259.020 211.800 ;
        RECT 260.720 3.300 262.320 211.800 ;
        RECT 264.020 3.300 265.620 211.800 ;
    END
  END vdda1
  PIN vssa1
    ANTENNADIFFAREA 167.107590 ;
    PORT
      LAYER pwell ;
        RECT 146.325 131.680 197.045 132.110 ;
        RECT 146.325 84.150 146.755 131.680 ;
        RECT 196.615 84.150 197.045 131.680 ;
        RECT 224.215 131.900 274.935 132.330 ;
        RECT 198.385 131.100 223.105 131.530 ;
        RECT 198.385 102.800 198.815 131.100 ;
        RECT 222.675 102.800 223.105 131.100 ;
        RECT 198.385 102.370 223.105 102.800 ;
        RECT 211.005 97.530 213.595 100.210 ;
        RECT 214.005 97.530 216.595 100.210 ;
        RECT 211.005 94.750 213.595 97.430 ;
        RECT 214.005 94.750 216.595 97.430 ;
        RECT 211.005 91.970 213.595 94.650 ;
        RECT 214.005 91.970 216.595 94.650 ;
        RECT 217.635 91.960 220.225 94.640 ;
        RECT 211.005 89.190 213.595 91.870 ;
        RECT 214.005 89.190 216.595 91.870 ;
        RECT 217.635 89.180 220.225 91.860 ;
        RECT 198.850 87.435 200.580 89.165 ;
        RECT 146.325 83.720 197.045 84.150 ;
        RECT 198.145 86.155 201.255 86.585 ;
        RECT 211.005 86.410 213.595 89.090 ;
        RECT 214.005 86.410 216.595 89.090 ;
        RECT 217.635 86.400 220.225 89.080 ;
        RECT 198.145 83.905 198.575 86.155 ;
        RECT 200.825 83.905 201.255 86.155 ;
        RECT 198.145 83.475 201.255 83.905 ;
        RECT 211.005 83.630 213.595 86.310 ;
        RECT 214.005 83.630 216.595 86.310 ;
        RECT 217.635 83.620 220.225 86.300 ;
        RECT 146.375 82.200 197.095 82.630 ;
        RECT 146.375 66.210 146.805 82.200 ;
        RECT 196.665 66.210 197.095 82.200 ;
        RECT 200.240 77.440 203.140 80.120 ;
        RECT 218.440 77.440 221.340 80.120 ;
        RECT 200.230 74.410 203.130 77.090 ;
        RECT 218.450 74.410 221.350 77.090 ;
        RECT 146.375 65.780 197.095 66.210 ;
        RECT 224.215 66.110 224.645 131.900 ;
        RECT 274.505 66.110 274.935 131.900 ;
        RECT 224.215 65.680 274.935 66.110 ;
      LAYER li1 ;
        RECT 228.355 132.200 248.235 132.260 ;
        RECT 224.345 132.030 274.805 132.200 ;
        RECT 151.145 131.980 170.960 131.985 ;
        RECT 146.455 131.810 196.915 131.980 ;
        RECT 146.455 84.020 146.625 131.810 ;
        RECT 196.745 89.030 196.915 131.810 ;
        RECT 199.625 131.400 220.285 131.565 ;
        RECT 198.515 131.230 222.975 131.400 ;
        RECT 198.515 102.670 198.685 131.230 ;
        RECT 199.625 131.200 220.285 131.230 ;
        RECT 222.805 102.670 222.975 131.230 ;
        RECT 198.515 102.500 222.975 102.670 ;
        RECT 210.695 100.020 211.290 100.045 ;
        RECT 213.260 100.020 214.250 100.050 ;
        RECT 216.265 100.020 217.950 100.075 ;
        RECT 210.695 99.850 217.950 100.020 ;
        RECT 210.695 97.890 211.365 99.850 ;
        RECT 213.235 97.890 214.365 99.850 ;
        RECT 214.915 98.390 215.375 98.560 ;
        RECT 216.235 97.890 217.950 99.850 ;
        RECT 210.695 97.070 217.950 97.890 ;
        RECT 210.695 95.110 211.365 97.070 ;
        RECT 213.235 95.110 214.365 97.070 ;
        RECT 214.915 95.610 215.375 95.780 ;
        RECT 216.235 95.110 217.950 97.070 ;
        RECT 210.695 94.450 217.950 95.110 ;
        RECT 210.695 94.290 220.035 94.450 ;
        RECT 210.695 92.330 211.365 94.290 ;
        RECT 213.235 92.330 214.365 94.290 ;
        RECT 216.235 94.280 220.035 94.290 ;
        RECT 214.915 92.830 215.375 93.000 ;
        RECT 216.235 92.330 217.995 94.280 ;
        RECT 218.545 92.820 219.005 92.990 ;
        RECT 210.695 92.320 217.995 92.330 ;
        RECT 219.865 92.320 220.035 94.280 ;
        RECT 210.695 91.510 220.035 92.320 ;
        RECT 210.695 89.550 211.365 91.510 ;
        RECT 213.235 89.550 214.365 91.510 ;
        RECT 216.235 91.500 220.035 91.510 ;
        RECT 214.915 90.050 215.375 90.220 ;
        RECT 216.235 89.550 217.995 91.500 ;
        RECT 218.545 90.830 219.005 91.000 ;
        RECT 210.695 89.540 217.995 89.550 ;
        RECT 219.865 89.540 220.035 91.500 ;
        RECT 210.695 89.370 220.035 89.540 ;
        RECT 198.980 89.030 200.450 89.035 ;
        RECT 196.745 88.865 200.760 89.030 ;
        RECT 196.745 87.735 199.150 88.865 ;
        RECT 200.270 87.735 200.760 88.865 ;
        RECT 196.745 87.670 200.760 87.735 ;
        RECT 210.695 88.890 220.020 89.370 ;
        RECT 210.695 88.730 220.035 88.890 ;
        RECT 196.745 87.115 200.765 87.670 ;
        RECT 196.745 86.285 201.285 87.115 ;
        RECT 151.240 84.020 171.055 84.060 ;
        RECT 196.745 84.020 198.445 86.285 ;
        RECT 146.455 83.850 198.445 84.020 ;
        RECT 151.240 83.800 171.055 83.850 ;
        RECT 198.275 83.775 198.445 83.850 ;
        RECT 200.945 83.775 201.285 86.285 ;
        RECT 210.695 86.770 211.365 88.730 ;
        RECT 213.235 86.770 214.365 88.730 ;
        RECT 216.235 88.720 220.035 88.730 ;
        RECT 214.915 87.270 215.375 87.440 ;
        RECT 216.235 86.770 217.995 88.720 ;
        RECT 218.545 87.260 219.005 87.430 ;
        RECT 210.695 86.760 217.995 86.770 ;
        RECT 219.865 86.760 220.035 88.720 ;
        RECT 210.695 86.590 220.035 86.760 ;
        RECT 210.695 86.110 220.020 86.590 ;
        RECT 210.695 85.950 220.035 86.110 ;
        RECT 210.695 83.990 211.365 85.950 ;
        RECT 213.235 83.990 214.365 85.950 ;
        RECT 216.235 85.940 220.035 85.950 ;
        RECT 214.915 84.490 215.375 84.660 ;
        RECT 216.235 83.990 217.995 85.940 ;
        RECT 210.695 83.980 217.995 83.990 ;
        RECT 219.865 83.980 220.035 85.940 ;
        RECT 210.695 83.845 220.035 83.980 ;
        RECT 210.695 83.840 213.405 83.845 ;
        RECT 211.195 83.820 213.405 83.840 ;
        RECT 214.195 83.830 220.035 83.845 ;
        RECT 214.195 83.820 216.405 83.830 ;
        RECT 217.825 83.810 220.035 83.830 ;
        RECT 198.275 83.605 201.285 83.775 ;
        RECT 151.240 82.500 171.055 82.545 ;
        RECT 146.505 82.330 196.965 82.500 ;
        RECT 146.505 66.080 146.675 82.330 ;
        RECT 151.240 82.285 171.055 82.330 ;
        RECT 151.215 66.080 171.030 66.120 ;
        RECT 196.795 66.080 196.965 82.330 ;
        RECT 199.790 79.740 203.280 80.370 ;
        RECT 199.790 77.810 200.620 79.740 ;
        RECT 201.460 79.090 201.920 79.260 ;
        RECT 202.750 77.810 203.280 79.740 ;
        RECT 199.790 76.730 203.280 77.810 ;
        RECT 199.790 74.790 200.620 76.730 ;
        RECT 201.450 75.270 201.910 75.440 ;
        RECT 202.750 74.790 203.280 76.730 ;
        RECT 199.790 74.160 203.280 74.790 ;
        RECT 218.300 79.740 221.790 80.370 ;
        RECT 218.300 77.810 218.830 79.740 ;
        RECT 219.660 79.090 220.120 79.260 ;
        RECT 220.960 77.810 221.790 79.740 ;
        RECT 218.300 76.730 221.790 77.810 ;
        RECT 218.300 74.790 218.830 76.730 ;
        RECT 219.670 75.270 220.130 75.440 ;
        RECT 220.960 74.790 221.790 76.730 ;
        RECT 218.300 74.160 221.790 74.790 ;
        RECT 146.505 65.910 196.965 66.080 ;
        RECT 224.345 65.980 224.515 132.030 ;
        RECT 228.355 132.000 248.235 132.030 ;
        RECT 228.365 65.980 248.245 66.030 ;
        RECT 274.635 65.980 274.805 132.030 ;
        RECT 151.215 65.860 171.030 65.910 ;
        RECT 224.345 65.810 274.805 65.980 ;
        RECT 228.365 65.770 248.245 65.810 ;
      LAYER mcon ;
        RECT 228.490 132.045 228.660 132.215 ;
        RECT 228.850 132.045 229.020 132.215 ;
        RECT 229.210 132.045 229.380 132.215 ;
        RECT 229.570 132.045 229.740 132.215 ;
        RECT 229.930 132.045 230.100 132.215 ;
        RECT 230.290 132.045 230.460 132.215 ;
        RECT 230.650 132.045 230.820 132.215 ;
        RECT 231.010 132.045 231.180 132.215 ;
        RECT 231.370 132.045 231.540 132.215 ;
        RECT 231.730 132.045 231.900 132.215 ;
        RECT 232.090 132.045 232.260 132.215 ;
        RECT 232.450 132.045 232.620 132.215 ;
        RECT 232.810 132.045 232.980 132.215 ;
        RECT 233.170 132.045 233.340 132.215 ;
        RECT 233.530 132.045 233.700 132.215 ;
        RECT 233.890 132.045 234.060 132.215 ;
        RECT 234.250 132.045 234.420 132.215 ;
        RECT 234.610 132.045 234.780 132.215 ;
        RECT 234.970 132.045 235.140 132.215 ;
        RECT 235.330 132.045 235.500 132.215 ;
        RECT 235.690 132.045 235.860 132.215 ;
        RECT 236.050 132.045 236.220 132.215 ;
        RECT 236.410 132.045 236.580 132.215 ;
        RECT 236.770 132.045 236.940 132.215 ;
        RECT 237.130 132.045 237.300 132.215 ;
        RECT 237.490 132.045 237.660 132.215 ;
        RECT 237.850 132.045 238.020 132.215 ;
        RECT 238.210 132.045 238.380 132.215 ;
        RECT 238.570 132.045 238.740 132.215 ;
        RECT 238.930 132.045 239.100 132.215 ;
        RECT 239.290 132.045 239.460 132.215 ;
        RECT 239.650 132.045 239.820 132.215 ;
        RECT 240.010 132.045 240.180 132.215 ;
        RECT 240.370 132.045 240.540 132.215 ;
        RECT 240.730 132.045 240.900 132.215 ;
        RECT 241.090 132.045 241.260 132.215 ;
        RECT 241.450 132.045 241.620 132.215 ;
        RECT 241.810 132.045 241.980 132.215 ;
        RECT 242.170 132.045 242.340 132.215 ;
        RECT 242.530 132.045 242.700 132.215 ;
        RECT 242.890 132.045 243.060 132.215 ;
        RECT 243.250 132.045 243.420 132.215 ;
        RECT 243.610 132.045 243.780 132.215 ;
        RECT 243.970 132.045 244.140 132.215 ;
        RECT 244.330 132.045 244.500 132.215 ;
        RECT 244.690 132.045 244.860 132.215 ;
        RECT 245.050 132.045 245.220 132.215 ;
        RECT 245.410 132.045 245.580 132.215 ;
        RECT 245.770 132.045 245.940 132.215 ;
        RECT 246.130 132.045 246.300 132.215 ;
        RECT 246.490 132.045 246.660 132.215 ;
        RECT 246.850 132.045 247.020 132.215 ;
        RECT 247.210 132.045 247.380 132.215 ;
        RECT 247.570 132.045 247.740 132.215 ;
        RECT 247.930 132.045 248.100 132.215 ;
        RECT 151.250 131.815 151.420 131.985 ;
        RECT 151.610 131.815 151.780 131.985 ;
        RECT 151.970 131.815 152.140 131.985 ;
        RECT 152.330 131.815 152.500 131.985 ;
        RECT 152.690 131.815 152.860 131.985 ;
        RECT 153.050 131.815 153.220 131.985 ;
        RECT 153.410 131.815 153.580 131.985 ;
        RECT 153.770 131.815 153.940 131.985 ;
        RECT 154.130 131.815 154.300 131.985 ;
        RECT 154.490 131.815 154.660 131.985 ;
        RECT 154.850 131.815 155.020 131.985 ;
        RECT 155.210 131.815 155.380 131.985 ;
        RECT 155.570 131.815 155.740 131.985 ;
        RECT 155.930 131.815 156.100 131.985 ;
        RECT 156.290 131.815 156.460 131.985 ;
        RECT 156.650 131.815 156.820 131.985 ;
        RECT 157.010 131.815 157.180 131.985 ;
        RECT 157.370 131.815 157.540 131.985 ;
        RECT 157.730 131.815 157.900 131.985 ;
        RECT 158.090 131.815 158.260 131.985 ;
        RECT 158.450 131.815 158.620 131.985 ;
        RECT 158.810 131.815 158.980 131.985 ;
        RECT 159.170 131.815 159.340 131.985 ;
        RECT 159.530 131.815 159.700 131.985 ;
        RECT 159.890 131.815 160.060 131.985 ;
        RECT 160.250 131.815 160.420 131.985 ;
        RECT 160.610 131.815 160.780 131.985 ;
        RECT 160.970 131.815 161.140 131.985 ;
        RECT 161.330 131.815 161.500 131.985 ;
        RECT 161.690 131.815 161.860 131.985 ;
        RECT 162.050 131.815 162.220 131.985 ;
        RECT 162.410 131.815 162.580 131.985 ;
        RECT 162.770 131.815 162.940 131.985 ;
        RECT 163.130 131.815 163.300 131.985 ;
        RECT 163.490 131.815 163.660 131.985 ;
        RECT 163.850 131.815 164.020 131.985 ;
        RECT 164.210 131.815 164.380 131.985 ;
        RECT 164.570 131.815 164.740 131.985 ;
        RECT 164.930 131.815 165.100 131.985 ;
        RECT 165.290 131.815 165.460 131.985 ;
        RECT 165.650 131.815 165.820 131.985 ;
        RECT 166.010 131.815 166.180 131.985 ;
        RECT 166.370 131.815 166.540 131.985 ;
        RECT 166.730 131.815 166.900 131.985 ;
        RECT 167.090 131.815 167.260 131.985 ;
        RECT 167.450 131.815 167.620 131.985 ;
        RECT 167.810 131.815 167.980 131.985 ;
        RECT 168.170 131.815 168.340 131.985 ;
        RECT 168.530 131.815 168.700 131.985 ;
        RECT 168.890 131.815 169.060 131.985 ;
        RECT 169.250 131.815 169.420 131.985 ;
        RECT 169.610 131.815 169.780 131.985 ;
        RECT 169.970 131.815 170.140 131.985 ;
        RECT 170.330 131.815 170.500 131.985 ;
        RECT 170.690 131.815 170.860 131.985 ;
        RECT 199.790 131.300 199.960 131.470 ;
        RECT 200.150 131.300 200.320 131.470 ;
        RECT 200.510 131.300 200.680 131.470 ;
        RECT 200.870 131.300 201.040 131.470 ;
        RECT 201.230 131.300 201.400 131.470 ;
        RECT 201.590 131.300 201.760 131.470 ;
        RECT 201.950 131.300 202.120 131.470 ;
        RECT 202.310 131.300 202.480 131.470 ;
        RECT 202.670 131.300 202.840 131.470 ;
        RECT 203.030 131.300 203.200 131.470 ;
        RECT 203.390 131.300 203.560 131.470 ;
        RECT 203.750 131.300 203.920 131.470 ;
        RECT 204.110 131.300 204.280 131.470 ;
        RECT 204.470 131.300 204.640 131.470 ;
        RECT 204.830 131.300 205.000 131.470 ;
        RECT 205.190 131.300 205.360 131.470 ;
        RECT 205.550 131.300 205.720 131.470 ;
        RECT 205.910 131.300 206.080 131.470 ;
        RECT 206.270 131.300 206.440 131.470 ;
        RECT 206.630 131.300 206.800 131.470 ;
        RECT 206.990 131.300 207.160 131.470 ;
        RECT 207.350 131.300 207.520 131.470 ;
        RECT 207.710 131.300 207.880 131.470 ;
        RECT 208.070 131.300 208.240 131.470 ;
        RECT 208.430 131.300 208.600 131.470 ;
        RECT 208.790 131.300 208.960 131.470 ;
        RECT 209.150 131.300 209.320 131.470 ;
        RECT 209.510 131.300 209.680 131.470 ;
        RECT 209.870 131.300 210.040 131.470 ;
        RECT 210.230 131.300 210.400 131.470 ;
        RECT 210.590 131.300 210.760 131.470 ;
        RECT 210.950 131.300 211.120 131.470 ;
        RECT 211.310 131.300 211.480 131.470 ;
        RECT 211.670 131.300 211.840 131.470 ;
        RECT 212.030 131.300 212.200 131.470 ;
        RECT 212.390 131.300 212.560 131.470 ;
        RECT 212.750 131.300 212.920 131.470 ;
        RECT 213.110 131.300 213.280 131.470 ;
        RECT 213.470 131.300 213.640 131.470 ;
        RECT 213.830 131.300 214.000 131.470 ;
        RECT 214.190 131.300 214.360 131.470 ;
        RECT 214.550 131.300 214.720 131.470 ;
        RECT 214.910 131.300 215.080 131.470 ;
        RECT 215.270 131.300 215.440 131.470 ;
        RECT 215.630 131.300 215.800 131.470 ;
        RECT 215.990 131.300 216.160 131.470 ;
        RECT 216.350 131.300 216.520 131.470 ;
        RECT 216.710 131.300 216.880 131.470 ;
        RECT 217.070 131.300 217.240 131.470 ;
        RECT 217.430 131.300 217.600 131.470 ;
        RECT 217.790 131.300 217.960 131.470 ;
        RECT 218.150 131.300 218.320 131.470 ;
        RECT 218.510 131.300 218.680 131.470 ;
        RECT 218.870 131.300 219.040 131.470 ;
        RECT 219.230 131.300 219.400 131.470 ;
        RECT 219.590 131.300 219.760 131.470 ;
        RECT 219.950 131.300 220.120 131.470 ;
        RECT 213.540 98.050 214.070 98.580 ;
        RECT 217.225 99.340 217.395 99.510 ;
        RECT 217.225 98.980 217.395 99.150 ;
        RECT 217.225 98.620 217.395 98.790 ;
        RECT 215.060 98.390 215.230 98.560 ;
        RECT 217.225 98.260 217.395 98.430 ;
        RECT 217.225 97.900 217.395 98.070 ;
        RECT 217.225 97.540 217.395 97.710 ;
        RECT 217.225 97.180 217.395 97.350 ;
        RECT 217.225 96.820 217.395 96.990 ;
        RECT 217.225 96.460 217.395 96.630 ;
        RECT 217.225 96.100 217.395 96.270 ;
        RECT 213.535 95.195 214.065 95.725 ;
        RECT 215.060 95.610 215.230 95.780 ;
        RECT 217.225 95.740 217.395 95.910 ;
        RECT 217.225 95.380 217.395 95.550 ;
        RECT 217.225 95.020 217.395 95.190 ;
        RECT 217.225 94.660 217.395 94.830 ;
        RECT 213.535 92.445 214.065 92.975 ;
        RECT 215.060 92.830 215.230 93.000 ;
        RECT 216.860 92.685 217.390 93.215 ;
        RECT 218.690 92.820 218.860 92.990 ;
        RECT 216.840 90.715 217.370 91.245 ;
        RECT 218.690 90.830 218.860 91.000 ;
        RECT 213.520 89.665 214.050 90.195 ;
        RECT 215.060 90.050 215.230 90.220 ;
        RECT 200.430 88.760 200.600 88.930 ;
        RECT 200.430 88.400 200.600 88.570 ;
        RECT 200.430 88.040 200.600 88.210 ;
        RECT 200.430 87.680 200.600 87.850 ;
        RECT 151.345 83.845 151.515 84.015 ;
        RECT 151.705 83.845 151.875 84.015 ;
        RECT 152.065 83.845 152.235 84.015 ;
        RECT 152.425 83.845 152.595 84.015 ;
        RECT 152.785 83.845 152.955 84.015 ;
        RECT 153.145 83.845 153.315 84.015 ;
        RECT 153.505 83.845 153.675 84.015 ;
        RECT 153.865 83.845 154.035 84.015 ;
        RECT 154.225 83.845 154.395 84.015 ;
        RECT 154.585 83.845 154.755 84.015 ;
        RECT 154.945 83.845 155.115 84.015 ;
        RECT 155.305 83.845 155.475 84.015 ;
        RECT 155.665 83.845 155.835 84.015 ;
        RECT 156.025 83.845 156.195 84.015 ;
        RECT 156.385 83.845 156.555 84.015 ;
        RECT 156.745 83.845 156.915 84.015 ;
        RECT 157.105 83.845 157.275 84.015 ;
        RECT 157.465 83.845 157.635 84.015 ;
        RECT 157.825 83.845 157.995 84.015 ;
        RECT 158.185 83.845 158.355 84.015 ;
        RECT 158.545 83.845 158.715 84.015 ;
        RECT 158.905 83.845 159.075 84.015 ;
        RECT 159.265 83.845 159.435 84.015 ;
        RECT 159.625 83.845 159.795 84.015 ;
        RECT 159.985 83.845 160.155 84.015 ;
        RECT 160.345 83.845 160.515 84.015 ;
        RECT 160.705 83.845 160.875 84.015 ;
        RECT 161.065 83.845 161.235 84.015 ;
        RECT 161.425 83.845 161.595 84.015 ;
        RECT 161.785 83.845 161.955 84.015 ;
        RECT 162.145 83.845 162.315 84.015 ;
        RECT 162.505 83.845 162.675 84.015 ;
        RECT 162.865 83.845 163.035 84.015 ;
        RECT 163.225 83.845 163.395 84.015 ;
        RECT 163.585 83.845 163.755 84.015 ;
        RECT 163.945 83.845 164.115 84.015 ;
        RECT 164.305 83.845 164.475 84.015 ;
        RECT 164.665 83.845 164.835 84.015 ;
        RECT 165.025 83.845 165.195 84.015 ;
        RECT 165.385 83.845 165.555 84.015 ;
        RECT 165.745 83.845 165.915 84.015 ;
        RECT 166.105 83.845 166.275 84.015 ;
        RECT 166.465 83.845 166.635 84.015 ;
        RECT 166.825 83.845 166.995 84.015 ;
        RECT 167.185 83.845 167.355 84.015 ;
        RECT 167.545 83.845 167.715 84.015 ;
        RECT 167.905 83.845 168.075 84.015 ;
        RECT 168.265 83.845 168.435 84.015 ;
        RECT 168.625 83.845 168.795 84.015 ;
        RECT 168.985 83.845 169.155 84.015 ;
        RECT 169.345 83.845 169.515 84.015 ;
        RECT 169.705 83.845 169.875 84.015 ;
        RECT 170.065 83.845 170.235 84.015 ;
        RECT 170.425 83.845 170.595 84.015 ;
        RECT 170.785 83.845 170.955 84.015 ;
        RECT 201.030 86.200 201.200 86.370 ;
        RECT 201.030 85.840 201.200 86.010 ;
        RECT 201.030 85.480 201.200 85.650 ;
        RECT 201.030 85.120 201.200 85.290 ;
        RECT 201.030 84.760 201.200 84.930 ;
        RECT 201.030 84.400 201.200 84.570 ;
        RECT 201.030 84.040 201.200 84.210 ;
        RECT 201.030 83.680 201.200 83.850 ;
        RECT 213.520 86.875 214.050 87.405 ;
        RECT 215.060 87.270 215.230 87.440 ;
        RECT 216.900 86.950 217.430 87.480 ;
        RECT 218.690 87.260 218.860 87.430 ;
        RECT 213.535 84.380 214.065 84.910 ;
        RECT 215.060 84.490 215.230 84.660 ;
        RECT 151.345 82.330 151.515 82.500 ;
        RECT 151.705 82.330 151.875 82.500 ;
        RECT 152.065 82.330 152.235 82.500 ;
        RECT 152.425 82.330 152.595 82.500 ;
        RECT 152.785 82.330 152.955 82.500 ;
        RECT 153.145 82.330 153.315 82.500 ;
        RECT 153.505 82.330 153.675 82.500 ;
        RECT 153.865 82.330 154.035 82.500 ;
        RECT 154.225 82.330 154.395 82.500 ;
        RECT 154.585 82.330 154.755 82.500 ;
        RECT 154.945 82.330 155.115 82.500 ;
        RECT 155.305 82.330 155.475 82.500 ;
        RECT 155.665 82.330 155.835 82.500 ;
        RECT 156.025 82.330 156.195 82.500 ;
        RECT 156.385 82.330 156.555 82.500 ;
        RECT 156.745 82.330 156.915 82.500 ;
        RECT 157.105 82.330 157.275 82.500 ;
        RECT 157.465 82.330 157.635 82.500 ;
        RECT 157.825 82.330 157.995 82.500 ;
        RECT 158.185 82.330 158.355 82.500 ;
        RECT 158.545 82.330 158.715 82.500 ;
        RECT 158.905 82.330 159.075 82.500 ;
        RECT 159.265 82.330 159.435 82.500 ;
        RECT 159.625 82.330 159.795 82.500 ;
        RECT 159.985 82.330 160.155 82.500 ;
        RECT 160.345 82.330 160.515 82.500 ;
        RECT 160.705 82.330 160.875 82.500 ;
        RECT 161.065 82.330 161.235 82.500 ;
        RECT 161.425 82.330 161.595 82.500 ;
        RECT 161.785 82.330 161.955 82.500 ;
        RECT 162.145 82.330 162.315 82.500 ;
        RECT 162.505 82.330 162.675 82.500 ;
        RECT 162.865 82.330 163.035 82.500 ;
        RECT 163.225 82.330 163.395 82.500 ;
        RECT 163.585 82.330 163.755 82.500 ;
        RECT 163.945 82.330 164.115 82.500 ;
        RECT 164.305 82.330 164.475 82.500 ;
        RECT 164.665 82.330 164.835 82.500 ;
        RECT 165.025 82.330 165.195 82.500 ;
        RECT 165.385 82.330 165.555 82.500 ;
        RECT 165.745 82.330 165.915 82.500 ;
        RECT 166.105 82.330 166.275 82.500 ;
        RECT 166.465 82.330 166.635 82.500 ;
        RECT 166.825 82.330 166.995 82.500 ;
        RECT 167.185 82.330 167.355 82.500 ;
        RECT 167.545 82.330 167.715 82.500 ;
        RECT 167.905 82.330 168.075 82.500 ;
        RECT 168.265 82.330 168.435 82.500 ;
        RECT 168.625 82.330 168.795 82.500 ;
        RECT 168.985 82.330 169.155 82.500 ;
        RECT 169.345 82.330 169.515 82.500 ;
        RECT 169.705 82.330 169.875 82.500 ;
        RECT 170.065 82.330 170.235 82.500 ;
        RECT 170.425 82.330 170.595 82.500 ;
        RECT 170.785 82.330 170.955 82.500 ;
        RECT 199.995 79.295 200.165 79.465 ;
        RECT 199.995 78.935 200.165 79.105 ;
        RECT 201.605 79.090 201.775 79.260 ;
        RECT 199.995 78.575 200.165 78.745 ;
        RECT 199.995 78.215 200.165 78.385 ;
        RECT 200.080 76.825 200.970 77.715 ;
        RECT 199.985 76.115 200.155 76.285 ;
        RECT 199.985 75.755 200.155 75.925 ;
        RECT 199.985 75.395 200.155 75.565 ;
        RECT 201.595 75.270 201.765 75.440 ;
        RECT 199.985 75.035 200.155 75.205 ;
        RECT 221.415 79.295 221.585 79.465 ;
        RECT 219.805 79.090 219.975 79.260 ;
        RECT 221.415 78.935 221.585 79.105 ;
        RECT 221.415 78.575 221.585 78.745 ;
        RECT 221.415 78.215 221.585 78.385 ;
        RECT 220.610 76.825 221.500 77.715 ;
        RECT 221.425 76.115 221.595 76.285 ;
        RECT 221.425 75.755 221.595 75.925 ;
        RECT 219.815 75.270 219.985 75.440 ;
        RECT 221.425 75.395 221.595 75.565 ;
        RECT 221.425 75.035 221.595 75.205 ;
        RECT 151.320 65.905 151.490 66.075 ;
        RECT 151.680 65.905 151.850 66.075 ;
        RECT 152.040 65.905 152.210 66.075 ;
        RECT 152.400 65.905 152.570 66.075 ;
        RECT 152.760 65.905 152.930 66.075 ;
        RECT 153.120 65.905 153.290 66.075 ;
        RECT 153.480 65.905 153.650 66.075 ;
        RECT 153.840 65.905 154.010 66.075 ;
        RECT 154.200 65.905 154.370 66.075 ;
        RECT 154.560 65.905 154.730 66.075 ;
        RECT 154.920 65.905 155.090 66.075 ;
        RECT 155.280 65.905 155.450 66.075 ;
        RECT 155.640 65.905 155.810 66.075 ;
        RECT 156.000 65.905 156.170 66.075 ;
        RECT 156.360 65.905 156.530 66.075 ;
        RECT 156.720 65.905 156.890 66.075 ;
        RECT 157.080 65.905 157.250 66.075 ;
        RECT 157.440 65.905 157.610 66.075 ;
        RECT 157.800 65.905 157.970 66.075 ;
        RECT 158.160 65.905 158.330 66.075 ;
        RECT 158.520 65.905 158.690 66.075 ;
        RECT 158.880 65.905 159.050 66.075 ;
        RECT 159.240 65.905 159.410 66.075 ;
        RECT 159.600 65.905 159.770 66.075 ;
        RECT 159.960 65.905 160.130 66.075 ;
        RECT 160.320 65.905 160.490 66.075 ;
        RECT 160.680 65.905 160.850 66.075 ;
        RECT 161.040 65.905 161.210 66.075 ;
        RECT 161.400 65.905 161.570 66.075 ;
        RECT 161.760 65.905 161.930 66.075 ;
        RECT 162.120 65.905 162.290 66.075 ;
        RECT 162.480 65.905 162.650 66.075 ;
        RECT 162.840 65.905 163.010 66.075 ;
        RECT 163.200 65.905 163.370 66.075 ;
        RECT 163.560 65.905 163.730 66.075 ;
        RECT 163.920 65.905 164.090 66.075 ;
        RECT 164.280 65.905 164.450 66.075 ;
        RECT 164.640 65.905 164.810 66.075 ;
        RECT 165.000 65.905 165.170 66.075 ;
        RECT 165.360 65.905 165.530 66.075 ;
        RECT 165.720 65.905 165.890 66.075 ;
        RECT 166.080 65.905 166.250 66.075 ;
        RECT 166.440 65.905 166.610 66.075 ;
        RECT 166.800 65.905 166.970 66.075 ;
        RECT 167.160 65.905 167.330 66.075 ;
        RECT 167.520 65.905 167.690 66.075 ;
        RECT 167.880 65.905 168.050 66.075 ;
        RECT 168.240 65.905 168.410 66.075 ;
        RECT 168.600 65.905 168.770 66.075 ;
        RECT 168.960 65.905 169.130 66.075 ;
        RECT 169.320 65.905 169.490 66.075 ;
        RECT 169.680 65.905 169.850 66.075 ;
        RECT 170.040 65.905 170.210 66.075 ;
        RECT 170.400 65.905 170.570 66.075 ;
        RECT 170.760 65.905 170.930 66.075 ;
        RECT 228.500 65.815 228.670 65.985 ;
        RECT 228.860 65.815 229.030 65.985 ;
        RECT 229.220 65.815 229.390 65.985 ;
        RECT 229.580 65.815 229.750 65.985 ;
        RECT 229.940 65.815 230.110 65.985 ;
        RECT 230.300 65.815 230.470 65.985 ;
        RECT 230.660 65.815 230.830 65.985 ;
        RECT 231.020 65.815 231.190 65.985 ;
        RECT 231.380 65.815 231.550 65.985 ;
        RECT 231.740 65.815 231.910 65.985 ;
        RECT 232.100 65.815 232.270 65.985 ;
        RECT 232.460 65.815 232.630 65.985 ;
        RECT 232.820 65.815 232.990 65.985 ;
        RECT 233.180 65.815 233.350 65.985 ;
        RECT 233.540 65.815 233.710 65.985 ;
        RECT 233.900 65.815 234.070 65.985 ;
        RECT 234.260 65.815 234.430 65.985 ;
        RECT 234.620 65.815 234.790 65.985 ;
        RECT 234.980 65.815 235.150 65.985 ;
        RECT 235.340 65.815 235.510 65.985 ;
        RECT 235.700 65.815 235.870 65.985 ;
        RECT 236.060 65.815 236.230 65.985 ;
        RECT 236.420 65.815 236.590 65.985 ;
        RECT 236.780 65.815 236.950 65.985 ;
        RECT 237.140 65.815 237.310 65.985 ;
        RECT 237.500 65.815 237.670 65.985 ;
        RECT 237.860 65.815 238.030 65.985 ;
        RECT 238.220 65.815 238.390 65.985 ;
        RECT 238.580 65.815 238.750 65.985 ;
        RECT 238.940 65.815 239.110 65.985 ;
        RECT 239.300 65.815 239.470 65.985 ;
        RECT 239.660 65.815 239.830 65.985 ;
        RECT 240.020 65.815 240.190 65.985 ;
        RECT 240.380 65.815 240.550 65.985 ;
        RECT 240.740 65.815 240.910 65.985 ;
        RECT 241.100 65.815 241.270 65.985 ;
        RECT 241.460 65.815 241.630 65.985 ;
        RECT 241.820 65.815 241.990 65.985 ;
        RECT 242.180 65.815 242.350 65.985 ;
        RECT 242.540 65.815 242.710 65.985 ;
        RECT 242.900 65.815 243.070 65.985 ;
        RECT 243.260 65.815 243.430 65.985 ;
        RECT 243.620 65.815 243.790 65.985 ;
        RECT 243.980 65.815 244.150 65.985 ;
        RECT 244.340 65.815 244.510 65.985 ;
        RECT 244.700 65.815 244.870 65.985 ;
        RECT 245.060 65.815 245.230 65.985 ;
        RECT 245.420 65.815 245.590 65.985 ;
        RECT 245.780 65.815 245.950 65.985 ;
        RECT 246.140 65.815 246.310 65.985 ;
        RECT 246.500 65.815 246.670 65.985 ;
        RECT 246.860 65.815 247.030 65.985 ;
        RECT 247.220 65.815 247.390 65.985 ;
        RECT 247.580 65.815 247.750 65.985 ;
        RECT 247.940 65.815 248.110 65.985 ;
      LAYER met1 ;
        RECT 228.355 132.290 248.235 132.310 ;
        RECT 151.145 132.015 170.960 132.075 ;
        RECT 151.085 131.780 171.020 132.015 ;
        RECT 228.295 131.970 248.295 132.290 ;
        RECT 228.355 131.950 248.235 131.970 ;
        RECT 151.145 131.715 170.960 131.780 ;
        RECT 199.625 131.595 220.285 131.615 ;
        RECT 199.565 131.170 220.345 131.595 ;
        RECT 199.625 131.150 220.285 131.170 ;
        RECT 213.320 98.445 214.290 98.760 ;
        RECT 214.935 98.445 215.355 98.590 ;
        RECT 213.320 98.360 215.355 98.445 ;
        RECT 213.320 98.185 215.345 98.360 ;
        RECT 213.320 97.870 214.290 98.185 ;
        RECT 213.315 95.625 214.285 95.905 ;
        RECT 214.935 95.625 215.355 95.810 ;
        RECT 213.315 95.365 215.355 95.625 ;
        RECT 213.315 95.015 214.285 95.365 ;
        RECT 217.020 94.475 217.600 99.690 ;
        RECT 216.700 93.395 217.550 93.415 ;
        RECT 213.315 92.855 214.285 93.155 ;
        RECT 214.935 92.855 215.355 93.030 ;
        RECT 216.640 92.860 217.610 93.395 ;
        RECT 218.565 92.860 218.985 93.020 ;
        RECT 213.315 92.595 215.365 92.855 ;
        RECT 216.640 92.600 219.010 92.860 ;
        RECT 213.315 92.265 214.285 92.595 ;
        RECT 216.640 92.505 217.610 92.600 ;
        RECT 216.700 92.485 217.550 92.505 ;
        RECT 216.680 91.425 217.530 91.445 ;
        RECT 216.620 91.195 217.590 91.425 ;
        RECT 216.620 90.935 219.000 91.195 ;
        RECT 216.620 90.535 217.590 90.935 ;
        RECT 218.565 90.800 218.985 90.935 ;
        RECT 216.680 90.515 217.530 90.535 ;
        RECT 213.300 90.085 214.270 90.375 ;
        RECT 214.935 90.085 215.355 90.250 ;
        RECT 213.300 89.825 215.375 90.085 ;
        RECT 213.300 89.485 214.270 89.825 ;
        RECT 200.240 88.985 200.790 89.090 ;
        RECT 200.240 87.680 202.925 88.985 ;
        RECT 200.240 87.520 200.790 87.680 ;
        RECT 200.915 86.050 201.315 86.505 ;
        RECT 201.835 86.050 202.920 87.680 ;
        RECT 216.740 87.660 217.590 87.680 ;
        RECT 213.300 87.280 214.270 87.585 ;
        RECT 214.935 87.280 215.355 87.470 ;
        RECT 213.300 87.240 215.355 87.280 ;
        RECT 216.680 87.370 217.650 87.660 ;
        RECT 218.565 87.370 218.985 87.460 ;
        RECT 213.300 87.020 215.330 87.240 ;
        RECT 216.680 87.110 218.990 87.370 ;
        RECT 213.300 86.695 214.270 87.020 ;
        RECT 216.680 86.770 217.650 87.110 ;
        RECT 216.740 86.750 217.590 86.770 ;
        RECT 200.915 84.265 202.920 86.050 ;
        RECT 213.315 84.535 214.285 85.090 ;
        RECT 214.935 84.535 215.355 84.690 ;
        RECT 200.915 84.180 202.925 84.265 ;
        RECT 213.315 84.235 215.365 84.535 ;
        RECT 213.315 84.200 214.285 84.235 ;
        RECT 151.240 84.090 171.055 84.110 ;
        RECT 151.180 83.770 171.115 84.090 ;
        RECT 151.240 83.750 171.055 83.770 ;
        RECT 200.915 83.545 201.315 84.180 ;
        RECT 201.835 83.825 202.925 84.180 ;
        RECT 151.240 82.575 171.055 82.595 ;
        RECT 151.180 82.255 171.115 82.575 ;
        RECT 151.240 82.235 171.055 82.255 ;
        RECT 208.770 81.565 209.760 81.585 ;
        RECT 198.650 79.580 199.650 81.505 ;
        RECT 208.745 80.595 212.890 81.565 ;
        RECT 208.770 80.575 209.760 80.595 ;
        RECT 211.885 80.565 212.845 80.595 ;
        RECT 221.930 79.580 222.930 81.505 ;
        RECT 198.650 79.160 201.910 79.580 ;
        RECT 219.670 79.160 222.930 79.580 ;
        RECT 198.650 78.050 200.740 79.160 ;
        RECT 201.480 79.060 201.900 79.160 ;
        RECT 219.680 79.060 220.100 79.160 ;
        RECT 220.840 78.050 222.930 79.160 ;
        RECT 198.650 76.500 201.110 78.050 ;
        RECT 220.470 76.500 222.930 78.050 ;
        RECT 198.650 75.340 200.740 76.500 ;
        RECT 201.470 75.340 201.890 75.470 ;
        RECT 219.690 75.340 220.110 75.470 ;
        RECT 220.840 75.340 222.930 76.500 ;
        RECT 198.650 74.920 201.900 75.340 ;
        RECT 219.680 74.920 222.930 75.340 ;
        RECT 198.650 74.065 199.650 74.920 ;
        RECT 221.930 74.065 222.930 74.920 ;
        RECT 151.215 66.150 171.030 66.170 ;
        RECT 151.155 65.830 171.090 66.150 ;
        RECT 228.365 66.060 248.245 66.080 ;
        RECT 151.215 65.810 171.030 65.830 ;
        RECT 228.305 65.740 248.305 66.060 ;
        RECT 228.365 65.720 248.245 65.740 ;
      LAYER via ;
        RECT 151.165 131.765 151.425 132.025 ;
        RECT 151.485 131.765 151.745 132.025 ;
        RECT 151.805 131.765 152.065 132.025 ;
        RECT 152.125 131.765 152.385 132.025 ;
        RECT 152.445 131.765 152.705 132.025 ;
        RECT 152.765 131.765 153.025 132.025 ;
        RECT 153.085 131.765 153.345 132.025 ;
        RECT 153.405 131.765 153.665 132.025 ;
        RECT 153.725 131.765 153.985 132.025 ;
        RECT 154.045 131.765 154.305 132.025 ;
        RECT 154.365 131.765 154.625 132.025 ;
        RECT 154.685 131.765 154.945 132.025 ;
        RECT 155.005 131.765 155.265 132.025 ;
        RECT 155.325 131.765 155.585 132.025 ;
        RECT 155.645 131.765 155.905 132.025 ;
        RECT 155.965 131.765 156.225 132.025 ;
        RECT 156.285 131.765 156.545 132.025 ;
        RECT 156.605 131.765 156.865 132.025 ;
        RECT 156.925 131.765 157.185 132.025 ;
        RECT 157.245 131.765 157.505 132.025 ;
        RECT 157.565 131.765 157.825 132.025 ;
        RECT 157.885 131.765 158.145 132.025 ;
        RECT 158.205 131.765 158.465 132.025 ;
        RECT 158.525 131.765 158.785 132.025 ;
        RECT 158.845 131.765 159.105 132.025 ;
        RECT 159.165 131.765 159.425 132.025 ;
        RECT 159.485 131.765 159.745 132.025 ;
        RECT 159.805 131.765 160.065 132.025 ;
        RECT 160.125 131.765 160.385 132.025 ;
        RECT 160.445 131.765 160.705 132.025 ;
        RECT 160.765 131.765 161.025 132.025 ;
        RECT 161.085 131.765 161.345 132.025 ;
        RECT 161.405 131.765 161.665 132.025 ;
        RECT 161.725 131.765 161.985 132.025 ;
        RECT 162.045 131.765 162.305 132.025 ;
        RECT 162.365 131.765 162.625 132.025 ;
        RECT 162.685 131.765 162.945 132.025 ;
        RECT 163.005 131.765 163.265 132.025 ;
        RECT 163.325 131.765 163.585 132.025 ;
        RECT 163.645 131.765 163.905 132.025 ;
        RECT 163.965 131.765 164.225 132.025 ;
        RECT 164.285 131.765 164.545 132.025 ;
        RECT 164.605 131.765 164.865 132.025 ;
        RECT 164.925 131.765 165.185 132.025 ;
        RECT 165.245 131.765 165.505 132.025 ;
        RECT 165.565 131.765 165.825 132.025 ;
        RECT 165.885 131.765 166.145 132.025 ;
        RECT 166.205 131.765 166.465 132.025 ;
        RECT 166.525 131.765 166.785 132.025 ;
        RECT 166.845 131.765 167.105 132.025 ;
        RECT 167.165 131.765 167.425 132.025 ;
        RECT 167.485 131.765 167.745 132.025 ;
        RECT 167.805 131.765 168.065 132.025 ;
        RECT 168.125 131.765 168.385 132.025 ;
        RECT 168.445 131.765 168.705 132.025 ;
        RECT 168.765 131.765 169.025 132.025 ;
        RECT 169.085 131.765 169.345 132.025 ;
        RECT 169.405 131.765 169.665 132.025 ;
        RECT 169.725 131.765 169.985 132.025 ;
        RECT 170.045 131.765 170.305 132.025 ;
        RECT 170.365 131.765 170.625 132.025 ;
        RECT 170.685 131.765 170.945 132.025 ;
        RECT 228.405 132.000 228.665 132.260 ;
        RECT 228.725 132.000 228.985 132.260 ;
        RECT 229.045 132.000 229.305 132.260 ;
        RECT 229.365 132.000 229.625 132.260 ;
        RECT 229.685 132.000 229.945 132.260 ;
        RECT 230.005 132.000 230.265 132.260 ;
        RECT 230.325 132.000 230.585 132.260 ;
        RECT 230.645 132.000 230.905 132.260 ;
        RECT 230.965 132.000 231.225 132.260 ;
        RECT 231.285 132.000 231.545 132.260 ;
        RECT 231.605 132.000 231.865 132.260 ;
        RECT 231.925 132.000 232.185 132.260 ;
        RECT 232.245 132.000 232.505 132.260 ;
        RECT 232.565 132.000 232.825 132.260 ;
        RECT 232.885 132.000 233.145 132.260 ;
        RECT 233.205 132.000 233.465 132.260 ;
        RECT 233.525 132.000 233.785 132.260 ;
        RECT 233.845 132.000 234.105 132.260 ;
        RECT 234.165 132.000 234.425 132.260 ;
        RECT 234.485 132.000 234.745 132.260 ;
        RECT 234.805 132.000 235.065 132.260 ;
        RECT 235.125 132.000 235.385 132.260 ;
        RECT 235.445 132.000 235.705 132.260 ;
        RECT 235.765 132.000 236.025 132.260 ;
        RECT 236.085 132.000 236.345 132.260 ;
        RECT 236.405 132.000 236.665 132.260 ;
        RECT 236.725 132.000 236.985 132.260 ;
        RECT 237.045 132.000 237.305 132.260 ;
        RECT 237.365 132.000 237.625 132.260 ;
        RECT 237.685 132.000 237.945 132.260 ;
        RECT 238.005 132.000 238.265 132.260 ;
        RECT 238.325 132.000 238.585 132.260 ;
        RECT 238.645 132.000 238.905 132.260 ;
        RECT 238.965 132.000 239.225 132.260 ;
        RECT 239.285 132.000 239.545 132.260 ;
        RECT 239.605 132.000 239.865 132.260 ;
        RECT 239.925 132.000 240.185 132.260 ;
        RECT 240.245 132.000 240.505 132.260 ;
        RECT 240.565 132.000 240.825 132.260 ;
        RECT 240.885 132.000 241.145 132.260 ;
        RECT 241.205 132.000 241.465 132.260 ;
        RECT 241.525 132.000 241.785 132.260 ;
        RECT 241.845 132.000 242.105 132.260 ;
        RECT 242.165 132.000 242.425 132.260 ;
        RECT 242.485 132.000 242.745 132.260 ;
        RECT 242.805 132.000 243.065 132.260 ;
        RECT 243.125 132.000 243.385 132.260 ;
        RECT 243.445 132.000 243.705 132.260 ;
        RECT 243.765 132.000 244.025 132.260 ;
        RECT 244.085 132.000 244.345 132.260 ;
        RECT 244.405 132.000 244.665 132.260 ;
        RECT 244.725 132.000 244.985 132.260 ;
        RECT 245.045 132.000 245.305 132.260 ;
        RECT 245.365 132.000 245.625 132.260 ;
        RECT 245.685 132.000 245.945 132.260 ;
        RECT 246.005 132.000 246.265 132.260 ;
        RECT 246.325 132.000 246.585 132.260 ;
        RECT 246.645 132.000 246.905 132.260 ;
        RECT 246.965 132.000 247.225 132.260 ;
        RECT 247.285 132.000 247.545 132.260 ;
        RECT 247.605 132.000 247.865 132.260 ;
        RECT 247.925 132.000 248.185 132.260 ;
        RECT 199.745 131.255 200.005 131.515 ;
        RECT 200.065 131.255 200.325 131.515 ;
        RECT 200.385 131.255 200.645 131.515 ;
        RECT 200.705 131.255 200.965 131.515 ;
        RECT 201.025 131.255 201.285 131.515 ;
        RECT 201.345 131.255 201.605 131.515 ;
        RECT 201.665 131.255 201.925 131.515 ;
        RECT 201.985 131.255 202.245 131.515 ;
        RECT 202.305 131.255 202.565 131.515 ;
        RECT 202.625 131.255 202.885 131.515 ;
        RECT 202.945 131.255 203.205 131.515 ;
        RECT 203.265 131.255 203.525 131.515 ;
        RECT 203.585 131.255 203.845 131.515 ;
        RECT 203.905 131.255 204.165 131.515 ;
        RECT 204.225 131.255 204.485 131.515 ;
        RECT 204.545 131.255 204.805 131.515 ;
        RECT 204.865 131.255 205.125 131.515 ;
        RECT 205.185 131.255 205.445 131.515 ;
        RECT 205.505 131.255 205.765 131.515 ;
        RECT 205.825 131.255 206.085 131.515 ;
        RECT 206.145 131.255 206.405 131.515 ;
        RECT 206.465 131.255 206.725 131.515 ;
        RECT 206.785 131.255 207.045 131.515 ;
        RECT 207.105 131.255 207.365 131.515 ;
        RECT 207.425 131.255 207.685 131.515 ;
        RECT 207.745 131.255 208.005 131.515 ;
        RECT 208.065 131.255 208.325 131.515 ;
        RECT 208.385 131.255 208.645 131.515 ;
        RECT 208.705 131.255 208.965 131.515 ;
        RECT 209.025 131.255 209.285 131.515 ;
        RECT 209.345 131.255 209.605 131.515 ;
        RECT 209.665 131.255 209.925 131.515 ;
        RECT 209.985 131.255 210.245 131.515 ;
        RECT 210.305 131.255 210.565 131.515 ;
        RECT 210.625 131.255 210.885 131.515 ;
        RECT 210.945 131.255 211.205 131.515 ;
        RECT 211.265 131.255 211.525 131.515 ;
        RECT 211.585 131.255 211.845 131.515 ;
        RECT 211.905 131.255 212.165 131.515 ;
        RECT 212.225 131.255 212.485 131.515 ;
        RECT 212.545 131.255 212.805 131.515 ;
        RECT 212.865 131.255 213.125 131.515 ;
        RECT 213.185 131.255 213.445 131.515 ;
        RECT 213.505 131.255 213.765 131.515 ;
        RECT 213.825 131.255 214.085 131.515 ;
        RECT 214.145 131.255 214.405 131.515 ;
        RECT 214.465 131.255 214.725 131.515 ;
        RECT 214.785 131.255 215.045 131.515 ;
        RECT 215.105 131.255 215.365 131.515 ;
        RECT 215.425 131.255 215.685 131.515 ;
        RECT 215.745 131.255 216.005 131.515 ;
        RECT 216.065 131.255 216.325 131.515 ;
        RECT 216.385 131.255 216.645 131.515 ;
        RECT 216.705 131.255 216.965 131.515 ;
        RECT 217.025 131.255 217.285 131.515 ;
        RECT 217.345 131.255 217.605 131.515 ;
        RECT 217.665 131.255 217.925 131.515 ;
        RECT 217.985 131.255 218.245 131.515 ;
        RECT 218.305 131.255 218.565 131.515 ;
        RECT 218.625 131.255 218.885 131.515 ;
        RECT 218.945 131.255 219.205 131.515 ;
        RECT 219.265 131.255 219.525 131.515 ;
        RECT 219.585 131.255 219.845 131.515 ;
        RECT 219.905 131.255 220.165 131.515 ;
        RECT 217.180 99.355 217.440 99.615 ;
        RECT 217.180 99.035 217.440 99.295 ;
        RECT 217.180 98.715 217.440 98.975 ;
        RECT 217.180 98.395 217.440 98.655 ;
        RECT 217.180 98.075 217.440 98.335 ;
        RECT 217.180 97.755 217.440 98.015 ;
        RECT 217.180 97.435 217.440 97.695 ;
        RECT 217.180 97.115 217.440 97.375 ;
        RECT 217.180 96.795 217.440 97.055 ;
        RECT 217.180 96.475 217.440 96.735 ;
        RECT 217.180 96.155 217.440 96.415 ;
        RECT 217.180 95.835 217.440 96.095 ;
        RECT 217.180 95.515 217.440 95.775 ;
        RECT 217.180 95.195 217.440 95.455 ;
        RECT 217.180 94.875 217.440 95.135 ;
        RECT 217.180 94.555 217.440 94.815 ;
        RECT 216.835 92.660 217.415 93.240 ;
        RECT 216.815 90.690 217.395 91.270 ;
        RECT 216.875 86.925 217.455 87.505 ;
        RECT 151.260 83.800 151.520 84.060 ;
        RECT 151.580 83.800 151.840 84.060 ;
        RECT 151.900 83.800 152.160 84.060 ;
        RECT 152.220 83.800 152.480 84.060 ;
        RECT 152.540 83.800 152.800 84.060 ;
        RECT 152.860 83.800 153.120 84.060 ;
        RECT 153.180 83.800 153.440 84.060 ;
        RECT 153.500 83.800 153.760 84.060 ;
        RECT 153.820 83.800 154.080 84.060 ;
        RECT 154.140 83.800 154.400 84.060 ;
        RECT 154.460 83.800 154.720 84.060 ;
        RECT 154.780 83.800 155.040 84.060 ;
        RECT 155.100 83.800 155.360 84.060 ;
        RECT 155.420 83.800 155.680 84.060 ;
        RECT 155.740 83.800 156.000 84.060 ;
        RECT 156.060 83.800 156.320 84.060 ;
        RECT 156.380 83.800 156.640 84.060 ;
        RECT 156.700 83.800 156.960 84.060 ;
        RECT 157.020 83.800 157.280 84.060 ;
        RECT 157.340 83.800 157.600 84.060 ;
        RECT 157.660 83.800 157.920 84.060 ;
        RECT 157.980 83.800 158.240 84.060 ;
        RECT 158.300 83.800 158.560 84.060 ;
        RECT 158.620 83.800 158.880 84.060 ;
        RECT 158.940 83.800 159.200 84.060 ;
        RECT 159.260 83.800 159.520 84.060 ;
        RECT 159.580 83.800 159.840 84.060 ;
        RECT 159.900 83.800 160.160 84.060 ;
        RECT 160.220 83.800 160.480 84.060 ;
        RECT 160.540 83.800 160.800 84.060 ;
        RECT 160.860 83.800 161.120 84.060 ;
        RECT 161.180 83.800 161.440 84.060 ;
        RECT 161.500 83.800 161.760 84.060 ;
        RECT 161.820 83.800 162.080 84.060 ;
        RECT 162.140 83.800 162.400 84.060 ;
        RECT 162.460 83.800 162.720 84.060 ;
        RECT 162.780 83.800 163.040 84.060 ;
        RECT 163.100 83.800 163.360 84.060 ;
        RECT 163.420 83.800 163.680 84.060 ;
        RECT 163.740 83.800 164.000 84.060 ;
        RECT 164.060 83.800 164.320 84.060 ;
        RECT 164.380 83.800 164.640 84.060 ;
        RECT 164.700 83.800 164.960 84.060 ;
        RECT 165.020 83.800 165.280 84.060 ;
        RECT 165.340 83.800 165.600 84.060 ;
        RECT 165.660 83.800 165.920 84.060 ;
        RECT 165.980 83.800 166.240 84.060 ;
        RECT 166.300 83.800 166.560 84.060 ;
        RECT 166.620 83.800 166.880 84.060 ;
        RECT 166.940 83.800 167.200 84.060 ;
        RECT 167.260 83.800 167.520 84.060 ;
        RECT 167.580 83.800 167.840 84.060 ;
        RECT 167.900 83.800 168.160 84.060 ;
        RECT 168.220 83.800 168.480 84.060 ;
        RECT 168.540 83.800 168.800 84.060 ;
        RECT 168.860 83.800 169.120 84.060 ;
        RECT 169.180 83.800 169.440 84.060 ;
        RECT 169.500 83.800 169.760 84.060 ;
        RECT 169.820 83.800 170.080 84.060 ;
        RECT 170.140 83.800 170.400 84.060 ;
        RECT 170.460 83.800 170.720 84.060 ;
        RECT 170.780 83.800 171.040 84.060 ;
        RECT 201.930 83.915 202.190 84.175 ;
        RECT 202.250 83.915 202.510 84.175 ;
        RECT 202.570 83.915 202.830 84.175 ;
        RECT 151.260 82.285 151.520 82.545 ;
        RECT 151.580 82.285 151.840 82.545 ;
        RECT 151.900 82.285 152.160 82.545 ;
        RECT 152.220 82.285 152.480 82.545 ;
        RECT 152.540 82.285 152.800 82.545 ;
        RECT 152.860 82.285 153.120 82.545 ;
        RECT 153.180 82.285 153.440 82.545 ;
        RECT 153.500 82.285 153.760 82.545 ;
        RECT 153.820 82.285 154.080 82.545 ;
        RECT 154.140 82.285 154.400 82.545 ;
        RECT 154.460 82.285 154.720 82.545 ;
        RECT 154.780 82.285 155.040 82.545 ;
        RECT 155.100 82.285 155.360 82.545 ;
        RECT 155.420 82.285 155.680 82.545 ;
        RECT 155.740 82.285 156.000 82.545 ;
        RECT 156.060 82.285 156.320 82.545 ;
        RECT 156.380 82.285 156.640 82.545 ;
        RECT 156.700 82.285 156.960 82.545 ;
        RECT 157.020 82.285 157.280 82.545 ;
        RECT 157.340 82.285 157.600 82.545 ;
        RECT 157.660 82.285 157.920 82.545 ;
        RECT 157.980 82.285 158.240 82.545 ;
        RECT 158.300 82.285 158.560 82.545 ;
        RECT 158.620 82.285 158.880 82.545 ;
        RECT 158.940 82.285 159.200 82.545 ;
        RECT 159.260 82.285 159.520 82.545 ;
        RECT 159.580 82.285 159.840 82.545 ;
        RECT 159.900 82.285 160.160 82.545 ;
        RECT 160.220 82.285 160.480 82.545 ;
        RECT 160.540 82.285 160.800 82.545 ;
        RECT 160.860 82.285 161.120 82.545 ;
        RECT 161.180 82.285 161.440 82.545 ;
        RECT 161.500 82.285 161.760 82.545 ;
        RECT 161.820 82.285 162.080 82.545 ;
        RECT 162.140 82.285 162.400 82.545 ;
        RECT 162.460 82.285 162.720 82.545 ;
        RECT 162.780 82.285 163.040 82.545 ;
        RECT 163.100 82.285 163.360 82.545 ;
        RECT 163.420 82.285 163.680 82.545 ;
        RECT 163.740 82.285 164.000 82.545 ;
        RECT 164.060 82.285 164.320 82.545 ;
        RECT 164.380 82.285 164.640 82.545 ;
        RECT 164.700 82.285 164.960 82.545 ;
        RECT 165.020 82.285 165.280 82.545 ;
        RECT 165.340 82.285 165.600 82.545 ;
        RECT 165.660 82.285 165.920 82.545 ;
        RECT 165.980 82.285 166.240 82.545 ;
        RECT 166.300 82.285 166.560 82.545 ;
        RECT 166.620 82.285 166.880 82.545 ;
        RECT 166.940 82.285 167.200 82.545 ;
        RECT 167.260 82.285 167.520 82.545 ;
        RECT 167.580 82.285 167.840 82.545 ;
        RECT 167.900 82.285 168.160 82.545 ;
        RECT 168.220 82.285 168.480 82.545 ;
        RECT 168.540 82.285 168.800 82.545 ;
        RECT 168.860 82.285 169.120 82.545 ;
        RECT 169.180 82.285 169.440 82.545 ;
        RECT 169.500 82.285 169.760 82.545 ;
        RECT 169.820 82.285 170.080 82.545 ;
        RECT 170.140 82.285 170.400 82.545 ;
        RECT 170.460 82.285 170.720 82.545 ;
        RECT 170.780 82.285 171.040 82.545 ;
        RECT 198.920 74.265 199.500 81.245 ;
        RECT 208.815 80.630 209.715 81.530 ;
        RECT 211.915 80.775 212.815 81.355 ;
        RECT 222.210 74.275 222.790 81.255 ;
        RECT 151.235 65.860 151.495 66.120 ;
        RECT 151.555 65.860 151.815 66.120 ;
        RECT 151.875 65.860 152.135 66.120 ;
        RECT 152.195 65.860 152.455 66.120 ;
        RECT 152.515 65.860 152.775 66.120 ;
        RECT 152.835 65.860 153.095 66.120 ;
        RECT 153.155 65.860 153.415 66.120 ;
        RECT 153.475 65.860 153.735 66.120 ;
        RECT 153.795 65.860 154.055 66.120 ;
        RECT 154.115 65.860 154.375 66.120 ;
        RECT 154.435 65.860 154.695 66.120 ;
        RECT 154.755 65.860 155.015 66.120 ;
        RECT 155.075 65.860 155.335 66.120 ;
        RECT 155.395 65.860 155.655 66.120 ;
        RECT 155.715 65.860 155.975 66.120 ;
        RECT 156.035 65.860 156.295 66.120 ;
        RECT 156.355 65.860 156.615 66.120 ;
        RECT 156.675 65.860 156.935 66.120 ;
        RECT 156.995 65.860 157.255 66.120 ;
        RECT 157.315 65.860 157.575 66.120 ;
        RECT 157.635 65.860 157.895 66.120 ;
        RECT 157.955 65.860 158.215 66.120 ;
        RECT 158.275 65.860 158.535 66.120 ;
        RECT 158.595 65.860 158.855 66.120 ;
        RECT 158.915 65.860 159.175 66.120 ;
        RECT 159.235 65.860 159.495 66.120 ;
        RECT 159.555 65.860 159.815 66.120 ;
        RECT 159.875 65.860 160.135 66.120 ;
        RECT 160.195 65.860 160.455 66.120 ;
        RECT 160.515 65.860 160.775 66.120 ;
        RECT 160.835 65.860 161.095 66.120 ;
        RECT 161.155 65.860 161.415 66.120 ;
        RECT 161.475 65.860 161.735 66.120 ;
        RECT 161.795 65.860 162.055 66.120 ;
        RECT 162.115 65.860 162.375 66.120 ;
        RECT 162.435 65.860 162.695 66.120 ;
        RECT 162.755 65.860 163.015 66.120 ;
        RECT 163.075 65.860 163.335 66.120 ;
        RECT 163.395 65.860 163.655 66.120 ;
        RECT 163.715 65.860 163.975 66.120 ;
        RECT 164.035 65.860 164.295 66.120 ;
        RECT 164.355 65.860 164.615 66.120 ;
        RECT 164.675 65.860 164.935 66.120 ;
        RECT 164.995 65.860 165.255 66.120 ;
        RECT 165.315 65.860 165.575 66.120 ;
        RECT 165.635 65.860 165.895 66.120 ;
        RECT 165.955 65.860 166.215 66.120 ;
        RECT 166.275 65.860 166.535 66.120 ;
        RECT 166.595 65.860 166.855 66.120 ;
        RECT 166.915 65.860 167.175 66.120 ;
        RECT 167.235 65.860 167.495 66.120 ;
        RECT 167.555 65.860 167.815 66.120 ;
        RECT 167.875 65.860 168.135 66.120 ;
        RECT 168.195 65.860 168.455 66.120 ;
        RECT 168.515 65.860 168.775 66.120 ;
        RECT 168.835 65.860 169.095 66.120 ;
        RECT 169.155 65.860 169.415 66.120 ;
        RECT 169.475 65.860 169.735 66.120 ;
        RECT 169.795 65.860 170.055 66.120 ;
        RECT 170.115 65.860 170.375 66.120 ;
        RECT 170.435 65.860 170.695 66.120 ;
        RECT 170.755 65.860 171.015 66.120 ;
        RECT 228.415 65.770 228.675 66.030 ;
        RECT 228.735 65.770 228.995 66.030 ;
        RECT 229.055 65.770 229.315 66.030 ;
        RECT 229.375 65.770 229.635 66.030 ;
        RECT 229.695 65.770 229.955 66.030 ;
        RECT 230.015 65.770 230.275 66.030 ;
        RECT 230.335 65.770 230.595 66.030 ;
        RECT 230.655 65.770 230.915 66.030 ;
        RECT 230.975 65.770 231.235 66.030 ;
        RECT 231.295 65.770 231.555 66.030 ;
        RECT 231.615 65.770 231.875 66.030 ;
        RECT 231.935 65.770 232.195 66.030 ;
        RECT 232.255 65.770 232.515 66.030 ;
        RECT 232.575 65.770 232.835 66.030 ;
        RECT 232.895 65.770 233.155 66.030 ;
        RECT 233.215 65.770 233.475 66.030 ;
        RECT 233.535 65.770 233.795 66.030 ;
        RECT 233.855 65.770 234.115 66.030 ;
        RECT 234.175 65.770 234.435 66.030 ;
        RECT 234.495 65.770 234.755 66.030 ;
        RECT 234.815 65.770 235.075 66.030 ;
        RECT 235.135 65.770 235.395 66.030 ;
        RECT 235.455 65.770 235.715 66.030 ;
        RECT 235.775 65.770 236.035 66.030 ;
        RECT 236.095 65.770 236.355 66.030 ;
        RECT 236.415 65.770 236.675 66.030 ;
        RECT 236.735 65.770 236.995 66.030 ;
        RECT 237.055 65.770 237.315 66.030 ;
        RECT 237.375 65.770 237.635 66.030 ;
        RECT 237.695 65.770 237.955 66.030 ;
        RECT 238.015 65.770 238.275 66.030 ;
        RECT 238.335 65.770 238.595 66.030 ;
        RECT 238.655 65.770 238.915 66.030 ;
        RECT 238.975 65.770 239.235 66.030 ;
        RECT 239.295 65.770 239.555 66.030 ;
        RECT 239.615 65.770 239.875 66.030 ;
        RECT 239.935 65.770 240.195 66.030 ;
        RECT 240.255 65.770 240.515 66.030 ;
        RECT 240.575 65.770 240.835 66.030 ;
        RECT 240.895 65.770 241.155 66.030 ;
        RECT 241.215 65.770 241.475 66.030 ;
        RECT 241.535 65.770 241.795 66.030 ;
        RECT 241.855 65.770 242.115 66.030 ;
        RECT 242.175 65.770 242.435 66.030 ;
        RECT 242.495 65.770 242.755 66.030 ;
        RECT 242.815 65.770 243.075 66.030 ;
        RECT 243.135 65.770 243.395 66.030 ;
        RECT 243.455 65.770 243.715 66.030 ;
        RECT 243.775 65.770 244.035 66.030 ;
        RECT 244.095 65.770 244.355 66.030 ;
        RECT 244.415 65.770 244.675 66.030 ;
        RECT 244.735 65.770 244.995 66.030 ;
        RECT 245.055 65.770 245.315 66.030 ;
        RECT 245.375 65.770 245.635 66.030 ;
        RECT 245.695 65.770 245.955 66.030 ;
        RECT 246.015 65.770 246.275 66.030 ;
        RECT 246.335 65.770 246.595 66.030 ;
        RECT 246.655 65.770 246.915 66.030 ;
        RECT 246.975 65.770 247.235 66.030 ;
        RECT 247.295 65.770 247.555 66.030 ;
        RECT 247.615 65.770 247.875 66.030 ;
        RECT 247.935 65.770 248.195 66.030 ;
      LAYER met2 ;
        RECT 151.100 132.025 171.100 134.100 ;
        RECT 151.095 131.765 171.100 132.025 ;
        RECT 228.285 131.985 248.285 134.100 ;
        RECT 151.100 84.060 171.100 131.765 ;
        RECT 198.985 130.965 248.285 131.985 ;
        RECT 201.930 103.085 219.490 130.965 ;
        RECT 228.285 100.815 248.285 130.965 ;
        RECT 216.515 94.785 248.285 100.815 ;
        RECT 216.515 90.260 221.645 94.785 ;
        RECT 218.880 89.950 221.645 90.260 ;
        RECT 228.285 89.950 248.285 94.785 ;
        RECT 218.880 88.535 248.285 89.950 ;
        RECT 216.530 86.555 248.285 88.535 ;
        RECT 151.100 83.800 171.105 84.060 ;
        RECT 201.785 83.875 202.975 84.215 ;
        RECT 222.310 83.920 248.285 86.555 ;
        RECT 151.100 82.545 171.100 83.800 ;
        RECT 151.100 82.285 171.105 82.545 ;
        RECT 151.100 63.930 171.100 82.285 ;
        RECT 201.835 81.530 202.920 83.875 ;
        RECT 208.720 81.530 209.810 81.535 ;
        RECT 196.635 80.625 209.810 81.530 ;
        RECT 211.835 81.475 212.895 81.510 ;
        RECT 228.285 81.475 248.285 83.920 ;
        RECT 196.635 80.550 209.765 80.625 ;
        RECT 211.835 80.615 248.285 81.475 ;
        RECT 211.880 80.590 248.285 80.615 ;
        RECT 196.635 74.075 199.665 80.550 ;
        RECT 221.910 74.050 248.285 80.590 ;
        RECT 228.285 66.030 248.285 74.050 ;
        RECT 228.285 65.770 248.295 66.030 ;
        RECT 228.285 63.930 248.285 65.770 ;
      LAYER via2 ;
        RECT 156.345 133.720 156.625 134.000 ;
        RECT 156.745 133.720 157.025 134.000 ;
        RECT 157.145 133.720 157.425 134.000 ;
        RECT 157.545 133.720 157.825 134.000 ;
        RECT 159.675 133.720 159.955 134.000 ;
        RECT 160.075 133.720 160.355 134.000 ;
        RECT 160.475 133.720 160.755 134.000 ;
        RECT 160.875 133.720 161.155 134.000 ;
        RECT 162.970 133.700 163.250 133.980 ;
        RECT 163.370 133.700 163.650 133.980 ;
        RECT 163.770 133.700 164.050 133.980 ;
        RECT 164.170 133.700 164.450 133.980 ;
        RECT 166.285 133.700 166.565 133.980 ;
        RECT 166.685 133.700 166.965 133.980 ;
        RECT 167.085 133.700 167.365 133.980 ;
        RECT 167.485 133.700 167.765 133.980 ;
        RECT 156.345 133.160 156.625 133.440 ;
        RECT 156.745 133.160 157.025 133.440 ;
        RECT 157.145 133.160 157.425 133.440 ;
        RECT 157.545 133.160 157.825 133.440 ;
        RECT 159.675 133.160 159.955 133.440 ;
        RECT 160.075 133.160 160.355 133.440 ;
        RECT 160.475 133.160 160.755 133.440 ;
        RECT 160.875 133.160 161.155 133.440 ;
        RECT 162.970 133.140 163.250 133.420 ;
        RECT 163.370 133.140 163.650 133.420 ;
        RECT 163.770 133.140 164.050 133.420 ;
        RECT 164.170 133.140 164.450 133.420 ;
        RECT 166.285 133.140 166.565 133.420 ;
        RECT 166.685 133.140 166.965 133.420 ;
        RECT 167.085 133.140 167.365 133.420 ;
        RECT 167.485 133.140 167.765 133.420 ;
        RECT 156.345 132.565 156.625 132.845 ;
        RECT 156.745 132.565 157.025 132.845 ;
        RECT 157.145 132.565 157.425 132.845 ;
        RECT 157.545 132.565 157.825 132.845 ;
        RECT 159.675 132.565 159.955 132.845 ;
        RECT 160.075 132.565 160.355 132.845 ;
        RECT 160.475 132.565 160.755 132.845 ;
        RECT 160.875 132.565 161.155 132.845 ;
        RECT 162.970 132.545 163.250 132.825 ;
        RECT 163.370 132.545 163.650 132.825 ;
        RECT 163.770 132.545 164.050 132.825 ;
        RECT 164.170 132.545 164.450 132.825 ;
        RECT 166.285 132.545 166.565 132.825 ;
        RECT 166.685 132.545 166.965 132.825 ;
        RECT 167.085 132.545 167.365 132.825 ;
        RECT 167.485 132.545 167.765 132.825 ;
        RECT 233.530 133.720 233.810 134.000 ;
        RECT 233.930 133.720 234.210 134.000 ;
        RECT 234.330 133.720 234.610 134.000 ;
        RECT 234.730 133.720 235.010 134.000 ;
        RECT 236.860 133.720 237.140 134.000 ;
        RECT 237.260 133.720 237.540 134.000 ;
        RECT 237.660 133.720 237.940 134.000 ;
        RECT 238.060 133.720 238.340 134.000 ;
        RECT 240.155 133.700 240.435 133.980 ;
        RECT 240.555 133.700 240.835 133.980 ;
        RECT 240.955 133.700 241.235 133.980 ;
        RECT 241.355 133.700 241.635 133.980 ;
        RECT 243.470 133.700 243.750 133.980 ;
        RECT 243.870 133.700 244.150 133.980 ;
        RECT 244.270 133.700 244.550 133.980 ;
        RECT 244.670 133.700 244.950 133.980 ;
        RECT 233.530 133.160 233.810 133.440 ;
        RECT 233.930 133.160 234.210 133.440 ;
        RECT 234.330 133.160 234.610 133.440 ;
        RECT 234.730 133.160 235.010 133.440 ;
        RECT 236.860 133.160 237.140 133.440 ;
        RECT 237.260 133.160 237.540 133.440 ;
        RECT 237.660 133.160 237.940 133.440 ;
        RECT 238.060 133.160 238.340 133.440 ;
        RECT 240.155 133.140 240.435 133.420 ;
        RECT 240.555 133.140 240.835 133.420 ;
        RECT 240.955 133.140 241.235 133.420 ;
        RECT 241.355 133.140 241.635 133.420 ;
        RECT 243.470 133.140 243.750 133.420 ;
        RECT 243.870 133.140 244.150 133.420 ;
        RECT 244.270 133.140 244.550 133.420 ;
        RECT 244.670 133.140 244.950 133.420 ;
        RECT 233.530 132.565 233.810 132.845 ;
        RECT 233.930 132.565 234.210 132.845 ;
        RECT 234.330 132.565 234.610 132.845 ;
        RECT 234.730 132.565 235.010 132.845 ;
        RECT 236.860 132.565 237.140 132.845 ;
        RECT 237.260 132.565 237.540 132.845 ;
        RECT 237.660 132.565 237.940 132.845 ;
        RECT 238.060 132.565 238.340 132.845 ;
        RECT 240.155 132.545 240.435 132.825 ;
        RECT 240.555 132.545 240.835 132.825 ;
        RECT 240.955 132.545 241.235 132.825 ;
        RECT 241.355 132.545 241.635 132.825 ;
        RECT 243.470 132.545 243.750 132.825 ;
        RECT 243.870 132.545 244.150 132.825 ;
        RECT 244.270 132.545 244.550 132.825 ;
        RECT 244.670 132.545 244.950 132.825 ;
        RECT 156.345 65.260 156.625 65.540 ;
        RECT 156.745 65.260 157.025 65.540 ;
        RECT 157.145 65.260 157.425 65.540 ;
        RECT 157.545 65.260 157.825 65.540 ;
        RECT 159.675 65.260 159.955 65.540 ;
        RECT 160.075 65.260 160.355 65.540 ;
        RECT 160.475 65.260 160.755 65.540 ;
        RECT 160.875 65.260 161.155 65.540 ;
        RECT 162.970 65.240 163.250 65.520 ;
        RECT 163.370 65.240 163.650 65.520 ;
        RECT 163.770 65.240 164.050 65.520 ;
        RECT 164.170 65.240 164.450 65.520 ;
        RECT 166.285 65.240 166.565 65.520 ;
        RECT 166.685 65.240 166.965 65.520 ;
        RECT 167.085 65.240 167.365 65.520 ;
        RECT 167.485 65.240 167.765 65.520 ;
        RECT 156.345 64.700 156.625 64.980 ;
        RECT 156.745 64.700 157.025 64.980 ;
        RECT 157.145 64.700 157.425 64.980 ;
        RECT 157.545 64.700 157.825 64.980 ;
        RECT 159.675 64.700 159.955 64.980 ;
        RECT 160.075 64.700 160.355 64.980 ;
        RECT 160.475 64.700 160.755 64.980 ;
        RECT 160.875 64.700 161.155 64.980 ;
        RECT 162.970 64.680 163.250 64.960 ;
        RECT 163.370 64.680 163.650 64.960 ;
        RECT 163.770 64.680 164.050 64.960 ;
        RECT 164.170 64.680 164.450 64.960 ;
        RECT 166.285 64.680 166.565 64.960 ;
        RECT 166.685 64.680 166.965 64.960 ;
        RECT 167.085 64.680 167.365 64.960 ;
        RECT 167.485 64.680 167.765 64.960 ;
        RECT 156.345 64.105 156.625 64.385 ;
        RECT 156.745 64.105 157.025 64.385 ;
        RECT 157.145 64.105 157.425 64.385 ;
        RECT 157.545 64.105 157.825 64.385 ;
        RECT 159.675 64.105 159.955 64.385 ;
        RECT 160.075 64.105 160.355 64.385 ;
        RECT 160.475 64.105 160.755 64.385 ;
        RECT 160.875 64.105 161.155 64.385 ;
        RECT 162.970 64.085 163.250 64.365 ;
        RECT 163.370 64.085 163.650 64.365 ;
        RECT 163.770 64.085 164.050 64.365 ;
        RECT 164.170 64.085 164.450 64.365 ;
        RECT 166.285 64.085 166.565 64.365 ;
        RECT 166.685 64.085 166.965 64.365 ;
        RECT 167.085 64.085 167.365 64.365 ;
        RECT 167.485 64.085 167.765 64.365 ;
        RECT 233.530 65.260 233.810 65.540 ;
        RECT 233.930 65.260 234.210 65.540 ;
        RECT 234.330 65.260 234.610 65.540 ;
        RECT 234.730 65.260 235.010 65.540 ;
        RECT 236.860 65.260 237.140 65.540 ;
        RECT 237.260 65.260 237.540 65.540 ;
        RECT 237.660 65.260 237.940 65.540 ;
        RECT 238.060 65.260 238.340 65.540 ;
        RECT 240.155 65.240 240.435 65.520 ;
        RECT 240.555 65.240 240.835 65.520 ;
        RECT 240.955 65.240 241.235 65.520 ;
        RECT 241.355 65.240 241.635 65.520 ;
        RECT 243.470 65.240 243.750 65.520 ;
        RECT 243.870 65.240 244.150 65.520 ;
        RECT 244.270 65.240 244.550 65.520 ;
        RECT 244.670 65.240 244.950 65.520 ;
        RECT 233.530 64.700 233.810 64.980 ;
        RECT 233.930 64.700 234.210 64.980 ;
        RECT 234.330 64.700 234.610 64.980 ;
        RECT 234.730 64.700 235.010 64.980 ;
        RECT 236.860 64.700 237.140 64.980 ;
        RECT 237.260 64.700 237.540 64.980 ;
        RECT 237.660 64.700 237.940 64.980 ;
        RECT 238.060 64.700 238.340 64.980 ;
        RECT 240.155 64.680 240.435 64.960 ;
        RECT 240.555 64.680 240.835 64.960 ;
        RECT 240.955 64.680 241.235 64.960 ;
        RECT 241.355 64.680 241.635 64.960 ;
        RECT 243.470 64.680 243.750 64.960 ;
        RECT 243.870 64.680 244.150 64.960 ;
        RECT 244.270 64.680 244.550 64.960 ;
        RECT 244.670 64.680 244.950 64.960 ;
        RECT 233.530 64.105 233.810 64.385 ;
        RECT 233.930 64.105 234.210 64.385 ;
        RECT 234.330 64.105 234.610 64.385 ;
        RECT 234.730 64.105 235.010 64.385 ;
        RECT 236.860 64.105 237.140 64.385 ;
        RECT 237.260 64.105 237.540 64.385 ;
        RECT 237.660 64.105 237.940 64.385 ;
        RECT 238.060 64.105 238.340 64.385 ;
        RECT 240.155 64.085 240.435 64.365 ;
        RECT 240.555 64.085 240.835 64.365 ;
        RECT 240.955 64.085 241.235 64.365 ;
        RECT 241.355 64.085 241.635 64.365 ;
        RECT 243.470 64.085 243.750 64.365 ;
        RECT 243.870 64.085 244.150 64.365 ;
        RECT 244.270 64.085 244.550 64.365 ;
        RECT 244.670 64.085 244.950 64.365 ;
      LAYER met3 ;
        RECT 151.100 132.390 171.100 134.100 ;
        RECT 228.285 132.390 248.285 134.100 ;
        RECT 151.100 63.930 171.100 65.640 ;
        RECT 228.285 63.930 248.285 65.640 ;
      LAYER via3 ;
        RECT 156.325 133.700 156.645 134.020 ;
        RECT 156.725 133.700 157.045 134.020 ;
        RECT 157.125 133.700 157.445 134.020 ;
        RECT 157.525 133.700 157.845 134.020 ;
        RECT 159.655 133.700 159.975 134.020 ;
        RECT 160.055 133.700 160.375 134.020 ;
        RECT 160.455 133.700 160.775 134.020 ;
        RECT 160.855 133.700 161.175 134.020 ;
        RECT 162.950 133.680 163.270 134.000 ;
        RECT 163.350 133.680 163.670 134.000 ;
        RECT 163.750 133.680 164.070 134.000 ;
        RECT 164.150 133.680 164.470 134.000 ;
        RECT 166.265 133.680 166.585 134.000 ;
        RECT 166.665 133.680 166.985 134.000 ;
        RECT 167.065 133.680 167.385 134.000 ;
        RECT 167.465 133.680 167.785 134.000 ;
        RECT 156.325 133.140 156.645 133.460 ;
        RECT 156.725 133.140 157.045 133.460 ;
        RECT 157.125 133.140 157.445 133.460 ;
        RECT 157.525 133.140 157.845 133.460 ;
        RECT 159.655 133.140 159.975 133.460 ;
        RECT 160.055 133.140 160.375 133.460 ;
        RECT 160.455 133.140 160.775 133.460 ;
        RECT 160.855 133.140 161.175 133.460 ;
        RECT 162.950 133.120 163.270 133.440 ;
        RECT 163.350 133.120 163.670 133.440 ;
        RECT 163.750 133.120 164.070 133.440 ;
        RECT 164.150 133.120 164.470 133.440 ;
        RECT 166.265 133.120 166.585 133.440 ;
        RECT 166.665 133.120 166.985 133.440 ;
        RECT 167.065 133.120 167.385 133.440 ;
        RECT 167.465 133.120 167.785 133.440 ;
        RECT 156.325 132.545 156.645 132.865 ;
        RECT 156.725 132.545 157.045 132.865 ;
        RECT 157.125 132.545 157.445 132.865 ;
        RECT 157.525 132.545 157.845 132.865 ;
        RECT 159.655 132.545 159.975 132.865 ;
        RECT 160.055 132.545 160.375 132.865 ;
        RECT 160.455 132.545 160.775 132.865 ;
        RECT 160.855 132.545 161.175 132.865 ;
        RECT 162.950 132.525 163.270 132.845 ;
        RECT 163.350 132.525 163.670 132.845 ;
        RECT 163.750 132.525 164.070 132.845 ;
        RECT 164.150 132.525 164.470 132.845 ;
        RECT 166.265 132.525 166.585 132.845 ;
        RECT 166.665 132.525 166.985 132.845 ;
        RECT 167.065 132.525 167.385 132.845 ;
        RECT 167.465 132.525 167.785 132.845 ;
        RECT 233.510 133.700 233.830 134.020 ;
        RECT 233.910 133.700 234.230 134.020 ;
        RECT 234.310 133.700 234.630 134.020 ;
        RECT 234.710 133.700 235.030 134.020 ;
        RECT 236.840 133.700 237.160 134.020 ;
        RECT 237.240 133.700 237.560 134.020 ;
        RECT 237.640 133.700 237.960 134.020 ;
        RECT 238.040 133.700 238.360 134.020 ;
        RECT 240.135 133.680 240.455 134.000 ;
        RECT 240.535 133.680 240.855 134.000 ;
        RECT 240.935 133.680 241.255 134.000 ;
        RECT 241.335 133.680 241.655 134.000 ;
        RECT 243.450 133.680 243.770 134.000 ;
        RECT 243.850 133.680 244.170 134.000 ;
        RECT 244.250 133.680 244.570 134.000 ;
        RECT 244.650 133.680 244.970 134.000 ;
        RECT 233.510 133.140 233.830 133.460 ;
        RECT 233.910 133.140 234.230 133.460 ;
        RECT 234.310 133.140 234.630 133.460 ;
        RECT 234.710 133.140 235.030 133.460 ;
        RECT 236.840 133.140 237.160 133.460 ;
        RECT 237.240 133.140 237.560 133.460 ;
        RECT 237.640 133.140 237.960 133.460 ;
        RECT 238.040 133.140 238.360 133.460 ;
        RECT 240.135 133.120 240.455 133.440 ;
        RECT 240.535 133.120 240.855 133.440 ;
        RECT 240.935 133.120 241.255 133.440 ;
        RECT 241.335 133.120 241.655 133.440 ;
        RECT 243.450 133.120 243.770 133.440 ;
        RECT 243.850 133.120 244.170 133.440 ;
        RECT 244.250 133.120 244.570 133.440 ;
        RECT 244.650 133.120 244.970 133.440 ;
        RECT 233.510 132.545 233.830 132.865 ;
        RECT 233.910 132.545 234.230 132.865 ;
        RECT 234.310 132.545 234.630 132.865 ;
        RECT 234.710 132.545 235.030 132.865 ;
        RECT 236.840 132.545 237.160 132.865 ;
        RECT 237.240 132.545 237.560 132.865 ;
        RECT 237.640 132.545 237.960 132.865 ;
        RECT 238.040 132.545 238.360 132.865 ;
        RECT 240.135 132.525 240.455 132.845 ;
        RECT 240.535 132.525 240.855 132.845 ;
        RECT 240.935 132.525 241.255 132.845 ;
        RECT 241.335 132.525 241.655 132.845 ;
        RECT 243.450 132.525 243.770 132.845 ;
        RECT 243.850 132.525 244.170 132.845 ;
        RECT 244.250 132.525 244.570 132.845 ;
        RECT 244.650 132.525 244.970 132.845 ;
        RECT 156.325 65.240 156.645 65.560 ;
        RECT 156.725 65.240 157.045 65.560 ;
        RECT 157.125 65.240 157.445 65.560 ;
        RECT 157.525 65.240 157.845 65.560 ;
        RECT 159.655 65.240 159.975 65.560 ;
        RECT 160.055 65.240 160.375 65.560 ;
        RECT 160.455 65.240 160.775 65.560 ;
        RECT 160.855 65.240 161.175 65.560 ;
        RECT 162.950 65.220 163.270 65.540 ;
        RECT 163.350 65.220 163.670 65.540 ;
        RECT 163.750 65.220 164.070 65.540 ;
        RECT 164.150 65.220 164.470 65.540 ;
        RECT 166.265 65.220 166.585 65.540 ;
        RECT 166.665 65.220 166.985 65.540 ;
        RECT 167.065 65.220 167.385 65.540 ;
        RECT 167.465 65.220 167.785 65.540 ;
        RECT 156.325 64.680 156.645 65.000 ;
        RECT 156.725 64.680 157.045 65.000 ;
        RECT 157.125 64.680 157.445 65.000 ;
        RECT 157.525 64.680 157.845 65.000 ;
        RECT 159.655 64.680 159.975 65.000 ;
        RECT 160.055 64.680 160.375 65.000 ;
        RECT 160.455 64.680 160.775 65.000 ;
        RECT 160.855 64.680 161.175 65.000 ;
        RECT 162.950 64.660 163.270 64.980 ;
        RECT 163.350 64.660 163.670 64.980 ;
        RECT 163.750 64.660 164.070 64.980 ;
        RECT 164.150 64.660 164.470 64.980 ;
        RECT 166.265 64.660 166.585 64.980 ;
        RECT 166.665 64.660 166.985 64.980 ;
        RECT 167.065 64.660 167.385 64.980 ;
        RECT 167.465 64.660 167.785 64.980 ;
        RECT 156.325 64.085 156.645 64.405 ;
        RECT 156.725 64.085 157.045 64.405 ;
        RECT 157.125 64.085 157.445 64.405 ;
        RECT 157.525 64.085 157.845 64.405 ;
        RECT 159.655 64.085 159.975 64.405 ;
        RECT 160.055 64.085 160.375 64.405 ;
        RECT 160.455 64.085 160.775 64.405 ;
        RECT 160.855 64.085 161.175 64.405 ;
        RECT 162.950 64.065 163.270 64.385 ;
        RECT 163.350 64.065 163.670 64.385 ;
        RECT 163.750 64.065 164.070 64.385 ;
        RECT 164.150 64.065 164.470 64.385 ;
        RECT 166.265 64.065 166.585 64.385 ;
        RECT 166.665 64.065 166.985 64.385 ;
        RECT 167.065 64.065 167.385 64.385 ;
        RECT 167.465 64.065 167.785 64.385 ;
        RECT 233.510 65.240 233.830 65.560 ;
        RECT 233.910 65.240 234.230 65.560 ;
        RECT 234.310 65.240 234.630 65.560 ;
        RECT 234.710 65.240 235.030 65.560 ;
        RECT 236.840 65.240 237.160 65.560 ;
        RECT 237.240 65.240 237.560 65.560 ;
        RECT 237.640 65.240 237.960 65.560 ;
        RECT 238.040 65.240 238.360 65.560 ;
        RECT 240.135 65.220 240.455 65.540 ;
        RECT 240.535 65.220 240.855 65.540 ;
        RECT 240.935 65.220 241.255 65.540 ;
        RECT 241.335 65.220 241.655 65.540 ;
        RECT 243.450 65.220 243.770 65.540 ;
        RECT 243.850 65.220 244.170 65.540 ;
        RECT 244.250 65.220 244.570 65.540 ;
        RECT 244.650 65.220 244.970 65.540 ;
        RECT 233.510 64.680 233.830 65.000 ;
        RECT 233.910 64.680 234.230 65.000 ;
        RECT 234.310 64.680 234.630 65.000 ;
        RECT 234.710 64.680 235.030 65.000 ;
        RECT 236.840 64.680 237.160 65.000 ;
        RECT 237.240 64.680 237.560 65.000 ;
        RECT 237.640 64.680 237.960 65.000 ;
        RECT 238.040 64.680 238.360 65.000 ;
        RECT 240.135 64.660 240.455 64.980 ;
        RECT 240.535 64.660 240.855 64.980 ;
        RECT 240.935 64.660 241.255 64.980 ;
        RECT 241.335 64.660 241.655 64.980 ;
        RECT 243.450 64.660 243.770 64.980 ;
        RECT 243.850 64.660 244.170 64.980 ;
        RECT 244.250 64.660 244.570 64.980 ;
        RECT 244.650 64.660 244.970 64.980 ;
        RECT 233.510 64.085 233.830 64.405 ;
        RECT 233.910 64.085 234.230 64.405 ;
        RECT 234.310 64.085 234.630 64.405 ;
        RECT 234.710 64.085 235.030 64.405 ;
        RECT 236.840 64.085 237.160 64.405 ;
        RECT 237.240 64.085 237.560 64.405 ;
        RECT 237.640 64.085 237.960 64.405 ;
        RECT 238.040 64.085 238.360 64.405 ;
        RECT 240.135 64.065 240.455 64.385 ;
        RECT 240.535 64.065 240.855 64.385 ;
        RECT 240.935 64.065 241.255 64.385 ;
        RECT 241.335 64.065 241.655 64.385 ;
        RECT 243.450 64.065 243.770 64.385 ;
        RECT 243.850 64.065 244.170 64.385 ;
        RECT 244.250 64.065 244.570 64.385 ;
        RECT 244.650 64.065 244.970 64.385 ;
      LAYER met4 ;
        RECT 156.315 3.300 157.915 211.800 ;
        RECT 159.615 3.300 161.215 211.800 ;
        RECT 162.915 3.300 164.515 211.800 ;
        RECT 166.215 3.300 167.815 211.800 ;
        RECT 233.500 3.300 235.100 211.800 ;
        RECT 236.800 3.300 238.400 211.800 ;
        RECT 240.100 3.300 241.700 211.800 ;
        RECT 243.400 3.300 245.000 211.800 ;
    END
  END vssa1
  PIN vssd1
    ANTENNADIFFAREA 15.428800 ;
    PORT
      LAYER pwell ;
        RECT 203.015 71.360 218.735 71.790 ;
        RECT 203.015 69.970 203.445 71.360 ;
        RECT 218.305 69.970 218.735 71.360 ;
        RECT 219.655 70.460 221.385 72.190 ;
        RECT 203.015 69.540 218.735 69.970 ;
        RECT 200.480 67.250 201.210 68.580 ;
        RECT 202.110 66.470 204.800 68.480 ;
        RECT 209.015 66.045 211.205 68.055 ;
        RECT 216.780 66.470 219.470 68.480 ;
        RECT 220.370 67.250 221.100 68.580 ;
        RECT 202.280 64.310 204.010 66.040 ;
        RECT 209.015 63.980 211.205 65.990 ;
        RECT 211.305 63.980 213.415 65.990 ;
      LAYER li1 ;
        RECT 219.785 71.890 221.255 72.060 ;
        RECT 203.145 71.490 218.605 71.660 ;
        RECT 203.145 69.840 203.315 71.490 ;
        RECT 218.435 69.840 218.605 71.490 ;
        RECT 203.145 69.670 218.605 69.840 ;
        RECT 219.785 70.760 219.955 71.890 ;
        RECT 221.085 70.760 221.255 71.890 ;
        RECT 219.785 70.590 221.255 70.760 ;
        RECT 203.145 69.140 218.595 69.670 ;
        RECT 219.785 68.980 220.800 70.590 ;
        RECT 201.920 68.410 204.670 68.560 ;
        RECT 200.610 68.180 204.670 68.410 ;
        RECT 200.610 67.060 202.430 68.180 ;
        RECT 202.780 67.170 203.820 67.340 ;
        RECT 201.920 66.770 202.430 67.060 ;
        RECT 204.500 66.770 204.670 68.180 ;
        RECT 216.910 68.410 219.660 68.560 ;
        RECT 216.910 68.180 220.970 68.410 ;
        RECT 211.080 67.925 211.430 67.930 ;
        RECT 201.920 66.600 204.670 66.770 ;
        RECT 209.145 67.755 211.445 67.925 ;
        RECT 201.920 66.570 203.875 66.600 ;
        RECT 201.960 65.910 203.875 66.570 ;
        RECT 209.145 66.345 209.315 67.755 ;
        RECT 209.995 67.185 210.535 67.355 ;
        RECT 210.905 66.345 211.445 67.755 ;
        RECT 216.910 66.770 217.080 68.180 ;
        RECT 217.760 67.170 218.800 67.340 ;
        RECT 219.150 67.060 220.970 68.180 ;
        RECT 219.150 66.770 219.660 67.060 ;
        RECT 216.910 66.600 219.660 66.770 ;
        RECT 219.150 66.570 219.660 66.600 ;
        RECT 209.145 66.175 211.445 66.345 ;
        RECT 201.960 65.740 203.880 65.910 ;
        RECT 209.150 65.860 211.445 66.175 ;
        RECT 201.960 64.610 202.580 65.740 ;
        RECT 203.710 64.610 203.880 65.740 ;
        RECT 201.960 64.445 203.880 64.610 ;
        RECT 202.410 64.440 203.880 64.445 ;
        RECT 209.145 65.690 213.285 65.860 ;
        RECT 209.145 64.280 209.315 65.690 ;
        RECT 210.905 64.280 211.605 65.690 ;
        RECT 212.285 65.120 212.745 65.290 ;
        RECT 213.115 64.280 213.285 65.690 ;
        RECT 209.145 64.110 213.285 64.280 ;
        RECT 211.070 64.060 211.445 64.110 ;
      LAYER mcon ;
        RECT 203.705 69.335 203.875 69.505 ;
        RECT 204.065 69.335 204.235 69.505 ;
        RECT 204.425 69.335 204.595 69.505 ;
        RECT 204.785 69.335 204.955 69.505 ;
        RECT 205.145 69.335 205.315 69.505 ;
        RECT 205.505 69.335 205.675 69.505 ;
        RECT 205.865 69.335 206.035 69.505 ;
        RECT 206.225 69.335 206.395 69.505 ;
        RECT 206.585 69.335 206.755 69.505 ;
        RECT 206.945 69.335 207.115 69.505 ;
        RECT 207.305 69.335 207.475 69.505 ;
        RECT 207.665 69.335 207.835 69.505 ;
        RECT 208.025 69.335 208.195 69.505 ;
        RECT 208.385 69.335 208.555 69.505 ;
        RECT 208.745 69.335 208.915 69.505 ;
        RECT 209.105 69.335 209.275 69.505 ;
        RECT 209.465 69.335 209.635 69.505 ;
        RECT 209.825 69.335 209.995 69.505 ;
        RECT 210.185 69.335 210.355 69.505 ;
        RECT 210.545 69.335 210.715 69.505 ;
        RECT 210.905 69.335 211.075 69.505 ;
        RECT 211.265 69.335 211.435 69.505 ;
        RECT 211.625 69.335 211.795 69.505 ;
        RECT 211.985 69.335 212.155 69.505 ;
        RECT 212.345 69.335 212.515 69.505 ;
        RECT 212.705 69.335 212.875 69.505 ;
        RECT 213.065 69.335 213.235 69.505 ;
        RECT 213.425 69.335 213.595 69.505 ;
        RECT 213.785 69.335 213.955 69.505 ;
        RECT 214.145 69.335 214.315 69.505 ;
        RECT 214.505 69.335 214.675 69.505 ;
        RECT 214.865 69.335 215.035 69.505 ;
        RECT 215.225 69.335 215.395 69.505 ;
        RECT 215.585 69.335 215.755 69.505 ;
        RECT 215.945 69.335 216.115 69.505 ;
        RECT 216.305 69.335 216.475 69.505 ;
        RECT 216.665 69.335 216.835 69.505 ;
        RECT 217.025 69.335 217.195 69.505 ;
        RECT 217.385 69.335 217.555 69.505 ;
        RECT 217.745 69.335 217.915 69.505 ;
        RECT 219.850 69.180 220.740 69.710 ;
        RECT 201.420 67.370 201.950 67.900 ;
        RECT 203.035 67.170 203.205 67.340 ;
        RECT 203.395 67.170 203.565 67.340 ;
        RECT 211.175 67.635 211.345 67.805 ;
        RECT 210.180 67.185 210.350 67.355 ;
        RECT 211.175 67.275 211.345 67.445 ;
        RECT 211.175 66.915 211.345 67.085 ;
        RECT 211.175 66.555 211.345 66.725 ;
        RECT 219.630 67.370 220.160 67.900 ;
        RECT 218.015 67.170 218.185 67.340 ;
        RECT 218.375 67.170 218.545 67.340 ;
        RECT 211.175 66.195 211.345 66.365 ;
        RECT 211.175 65.835 211.345 66.005 ;
        RECT 211.175 65.475 211.345 65.645 ;
        RECT 211.175 65.115 211.345 65.285 ;
        RECT 212.430 65.120 212.600 65.290 ;
      LAYER met1 ;
        RECT 201.385 68.810 220.800 69.910 ;
        RECT 201.385 68.500 202.395 68.810 ;
        RECT 201.340 67.160 202.395 68.500 ;
        RECT 210.030 68.370 212.745 68.810 ;
        RECT 219.640 68.500 220.800 68.810 ;
        RECT 210.030 67.385 210.490 68.370 ;
        RECT 201.340 67.150 202.400 67.160 ;
        RECT 202.800 67.150 203.800 67.370 ;
        RECT 210.015 67.155 210.515 67.385 ;
        RECT 201.340 66.920 203.810 67.150 ;
        RECT 201.340 66.260 202.395 66.920 ;
        RECT 211.075 65.010 211.455 68.370 ;
        RECT 212.310 65.320 212.745 68.370 ;
        RECT 217.780 67.150 218.780 67.370 ;
        RECT 219.240 67.160 220.800 68.500 ;
        RECT 219.180 67.150 220.800 67.160 ;
        RECT 217.770 66.920 220.800 67.150 ;
        RECT 219.240 66.270 220.800 66.920 ;
        RECT 219.240 66.260 220.240 66.270 ;
        RECT 212.305 65.100 212.745 65.320 ;
        RECT 212.305 65.090 212.725 65.100 ;
      LAYER via ;
        RECT 201.610 66.490 202.190 67.070 ;
      LAYER met2 ;
        RECT 201.395 63.930 202.395 68.590 ;
      LAYER via2 ;
        RECT 201.595 67.820 201.875 68.100 ;
        RECT 201.995 67.820 202.275 68.100 ;
        RECT 201.595 67.225 201.875 67.505 ;
        RECT 201.995 67.225 202.275 67.505 ;
        RECT 201.595 66.620 201.875 66.900 ;
        RECT 201.995 66.620 202.275 66.900 ;
        RECT 201.595 66.085 201.875 66.365 ;
        RECT 201.995 66.085 202.275 66.365 ;
        RECT 201.595 65.455 201.875 65.735 ;
        RECT 201.995 65.455 202.275 65.735 ;
        RECT 201.595 64.895 201.875 65.175 ;
        RECT 201.995 64.895 202.275 65.175 ;
        RECT 201.595 64.300 201.875 64.580 ;
        RECT 201.995 64.300 202.275 64.580 ;
      LAYER met3 ;
        RECT 201.395 63.930 202.395 68.590 ;
      LAYER via3 ;
        RECT 201.575 67.800 201.895 68.120 ;
        RECT 201.975 67.800 202.295 68.120 ;
        RECT 201.575 67.205 201.895 67.525 ;
        RECT 201.975 67.205 202.295 67.525 ;
        RECT 201.575 66.600 201.895 66.920 ;
        RECT 201.975 66.600 202.295 66.920 ;
        RECT 201.575 66.065 201.895 66.385 ;
        RECT 201.975 66.065 202.295 66.385 ;
        RECT 201.575 65.435 201.895 65.755 ;
        RECT 201.975 65.435 202.295 65.755 ;
        RECT 201.575 64.875 201.895 65.195 ;
        RECT 201.975 64.875 202.295 65.195 ;
        RECT 201.575 64.280 201.895 64.600 ;
        RECT 201.975 64.280 202.295 64.600 ;
      LAYER met4 ;
        RECT 201.105 3.300 202.705 211.800 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER nwell ;
        RECT 204.890 66.420 207.730 68.530 ;
        RECT 213.850 66.420 216.690 68.530 ;
        RECT 204.935 63.930 207.775 66.420 ;
      LAYER li1 ;
        RECT 207.935 97.910 208.395 98.080 ;
        RECT 205.070 68.180 207.910 68.570 ;
        RECT 205.070 66.770 205.240 68.180 ;
        RECT 207.380 67.840 207.910 68.180 ;
        RECT 213.670 68.180 216.510 68.570 ;
        RECT 213.670 67.840 214.200 68.180 ;
        RECT 205.970 67.170 207.010 67.340 ;
        RECT 207.380 67.050 208.370 67.840 ;
        RECT 213.210 67.050 214.200 67.840 ;
        RECT 214.570 67.170 215.610 67.340 ;
        RECT 207.380 66.770 207.910 67.050 ;
        RECT 205.070 66.600 207.910 66.770 ;
        RECT 205.115 66.580 207.910 66.600 ;
        RECT 213.670 66.770 214.200 67.050 ;
        RECT 216.340 66.770 216.510 68.180 ;
        RECT 213.670 66.600 216.510 66.770 ;
        RECT 213.670 66.580 214.180 66.600 ;
        RECT 205.115 65.690 207.595 66.580 ;
        RECT 205.115 64.280 205.285 65.690 ;
        RECT 205.655 65.120 206.695 65.290 ;
        RECT 207.425 64.280 207.595 65.690 ;
        RECT 205.115 64.110 207.595 64.280 ;
      LAYER mcon ;
        RECT 208.080 97.910 208.250 98.080 ;
        RECT 206.225 67.170 206.395 67.340 ;
        RECT 206.585 67.170 206.755 67.340 ;
        RECT 207.700 67.200 208.230 67.730 ;
        RECT 213.350 67.200 213.880 67.730 ;
        RECT 214.825 67.170 214.995 67.340 ;
        RECT 215.185 67.170 215.355 67.340 ;
        RECT 205.910 65.120 206.080 65.290 ;
        RECT 206.270 65.120 206.440 65.290 ;
      LAYER met1 ;
        RECT 207.955 97.955 208.375 98.110 ;
        RECT 210.745 97.955 211.550 98.185 ;
        RECT 207.940 97.580 211.550 97.955 ;
        RECT 210.745 97.300 211.550 97.580 ;
        RECT 205.990 67.200 206.990 67.370 ;
        RECT 207.370 67.200 208.370 68.520 ;
        RECT 205.990 66.970 208.370 67.200 ;
        RECT 207.370 66.130 208.370 66.970 ;
        RECT 213.210 67.200 214.210 68.520 ;
        RECT 214.590 67.200 215.590 67.370 ;
        RECT 213.210 66.970 215.590 67.200 ;
        RECT 213.210 66.130 214.210 66.970 ;
        RECT 207.415 65.540 208.415 66.130 ;
        RECT 205.695 65.320 208.415 65.540 ;
        RECT 205.675 65.275 208.415 65.320 ;
        RECT 205.675 65.090 206.675 65.275 ;
      LAYER via ;
        RECT 210.860 97.455 211.440 98.035 ;
        RECT 207.620 67.365 208.200 68.265 ;
        RECT 213.475 66.340 214.055 66.920 ;
      LAYER met2 ;
        RECT 210.745 98.135 211.550 98.180 ;
        RECT 210.695 97.350 211.600 98.135 ;
        RECT 207.425 67.875 208.415 68.530 ;
        RECT 210.745 67.875 211.550 97.350 ;
        RECT 207.425 67.125 214.770 67.875 ;
        RECT 207.435 67.045 214.770 67.125 ;
        RECT 213.270 66.215 214.770 67.045 ;
        RECT 213.770 63.930 214.770 66.215 ;
      LAYER via2 ;
        RECT 213.970 67.540 214.250 67.820 ;
        RECT 214.370 67.540 214.650 67.820 ;
        RECT 213.970 66.925 214.250 67.205 ;
        RECT 214.370 66.925 214.650 67.205 ;
        RECT 213.970 66.365 214.250 66.645 ;
        RECT 214.370 66.365 214.650 66.645 ;
        RECT 213.970 65.770 214.250 66.050 ;
        RECT 214.370 65.770 214.650 66.050 ;
        RECT 213.970 65.150 214.250 65.430 ;
        RECT 214.370 65.150 214.650 65.430 ;
        RECT 213.970 64.615 214.250 64.895 ;
        RECT 214.370 64.615 214.650 64.895 ;
      LAYER met3 ;
        RECT 213.770 63.930 214.770 67.875 ;
      LAYER via3 ;
        RECT 213.950 67.520 214.270 67.840 ;
        RECT 214.350 67.520 214.670 67.840 ;
        RECT 213.950 66.905 214.270 67.225 ;
        RECT 214.350 66.905 214.670 67.225 ;
        RECT 213.950 66.345 214.270 66.665 ;
        RECT 214.350 66.345 214.670 66.665 ;
        RECT 213.950 65.750 214.270 66.070 ;
        RECT 214.350 65.750 214.670 66.070 ;
        RECT 213.950 65.130 214.270 65.450 ;
        RECT 214.350 65.130 214.670 65.450 ;
        RECT 213.950 64.595 214.270 64.915 ;
        RECT 214.350 64.595 214.670 64.915 ;
      LAYER met4 ;
        RECT 213.440 3.300 215.040 211.800 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 198.780 74.430 199.520 80.460 ;
        RECT 222.060 74.430 222.800 80.460 ;
      LAYER li1 ;
        RECT 147.105 130.980 149.265 131.330 ;
        RECT 194.105 130.980 196.265 131.330 ;
        RECT 224.995 131.200 227.155 131.550 ;
        RECT 147.105 130.150 149.265 130.500 ;
        RECT 194.105 130.150 196.265 130.500 ;
        RECT 199.165 130.060 201.325 130.750 ;
        RECT 224.995 130.370 227.155 130.720 ;
        RECT 271.995 130.370 274.155 130.720 ;
        RECT 147.105 129.320 149.265 129.670 ;
        RECT 194.105 129.320 196.265 129.670 ;
        RECT 199.165 128.890 201.325 129.580 ;
        RECT 220.165 128.890 222.325 129.580 ;
        RECT 224.995 129.540 227.155 129.890 ;
        RECT 271.995 129.540 274.155 129.890 ;
        RECT 147.105 128.490 149.265 128.840 ;
        RECT 194.105 128.490 196.265 128.840 ;
        RECT 224.995 128.710 227.155 129.060 ;
        RECT 271.995 128.710 274.155 129.060 ;
        RECT 147.105 127.660 149.265 128.010 ;
        RECT 194.105 127.660 196.265 128.010 ;
        RECT 199.165 127.720 201.325 128.410 ;
        RECT 220.165 127.720 222.325 128.410 ;
        RECT 224.995 127.880 227.155 128.230 ;
        RECT 271.995 127.880 274.155 128.230 ;
        RECT 147.105 126.830 149.265 127.180 ;
        RECT 194.105 126.830 196.265 127.180 ;
        RECT 199.165 126.550 201.325 127.240 ;
        RECT 220.165 126.550 222.325 127.240 ;
        RECT 224.995 127.050 227.155 127.400 ;
        RECT 271.995 127.050 274.155 127.400 ;
        RECT 147.105 126.000 149.265 126.350 ;
        RECT 194.105 126.000 196.265 126.350 ;
        RECT 224.995 126.220 227.155 126.570 ;
        RECT 271.995 126.220 274.155 126.570 ;
        RECT 147.105 125.170 149.265 125.520 ;
        RECT 194.105 125.170 196.265 125.520 ;
        RECT 199.165 125.380 201.325 126.070 ;
        RECT 220.165 125.380 222.325 126.070 ;
        RECT 224.995 125.390 227.155 125.740 ;
        RECT 271.995 125.390 274.155 125.740 ;
        RECT 147.105 124.340 149.265 124.690 ;
        RECT 194.105 124.340 196.265 124.690 ;
        RECT 199.165 124.210 201.325 124.900 ;
        RECT 220.165 124.210 222.325 124.900 ;
        RECT 224.995 124.560 227.155 124.910 ;
        RECT 271.995 124.560 274.155 124.910 ;
        RECT 147.105 123.510 149.265 123.860 ;
        RECT 194.105 123.510 196.265 123.860 ;
        RECT 224.995 123.730 227.155 124.080 ;
        RECT 271.995 123.730 274.155 124.080 ;
        RECT 199.165 123.040 201.325 123.730 ;
        RECT 220.165 123.040 222.325 123.730 ;
        RECT 147.105 122.680 149.265 123.030 ;
        RECT 194.105 122.680 196.265 123.030 ;
        RECT 224.995 122.900 227.155 123.250 ;
        RECT 271.995 122.900 274.155 123.250 ;
        RECT 147.105 121.850 149.265 122.200 ;
        RECT 194.105 121.850 196.265 122.200 ;
        RECT 199.165 121.870 201.325 122.560 ;
        RECT 220.165 121.870 222.325 122.560 ;
        RECT 224.995 122.070 227.155 122.420 ;
        RECT 271.995 122.070 274.155 122.420 ;
        RECT 147.105 121.020 149.265 121.370 ;
        RECT 194.105 121.020 196.265 121.370 ;
        RECT 199.165 120.700 201.325 121.390 ;
        RECT 220.165 120.700 222.325 121.390 ;
        RECT 224.995 121.240 227.155 121.590 ;
        RECT 271.995 121.240 274.155 121.590 ;
        RECT 147.105 120.190 149.265 120.540 ;
        RECT 194.105 120.190 196.265 120.540 ;
        RECT 224.995 120.410 227.155 120.760 ;
        RECT 271.995 120.410 274.155 120.760 ;
        RECT 147.105 119.360 149.265 119.710 ;
        RECT 194.105 119.360 196.265 119.710 ;
        RECT 199.165 119.530 201.325 120.220 ;
        RECT 220.165 119.530 222.325 120.220 ;
        RECT 224.995 119.580 227.155 119.930 ;
        RECT 271.995 119.580 274.155 119.930 ;
        RECT 147.105 118.530 149.265 118.880 ;
        RECT 194.105 118.530 196.265 118.880 ;
        RECT 199.165 118.360 201.325 119.050 ;
        RECT 220.165 118.360 222.325 119.050 ;
        RECT 224.995 118.750 227.155 119.100 ;
        RECT 271.995 118.750 274.155 119.100 ;
        RECT 147.105 117.700 149.265 118.050 ;
        RECT 194.105 117.700 196.265 118.050 ;
        RECT 224.995 117.920 227.155 118.270 ;
        RECT 271.995 117.920 274.155 118.270 ;
        RECT 147.105 116.870 149.265 117.220 ;
        RECT 194.105 116.870 196.265 117.220 ;
        RECT 199.165 117.190 201.325 117.880 ;
        RECT 220.165 117.190 222.325 117.880 ;
        RECT 224.995 117.090 227.155 117.440 ;
        RECT 271.995 117.090 274.155 117.440 ;
        RECT 147.105 116.040 149.265 116.390 ;
        RECT 194.105 116.040 196.265 116.390 ;
        RECT 199.165 116.020 201.325 116.710 ;
        RECT 220.165 116.020 222.325 116.710 ;
        RECT 224.995 116.260 227.155 116.610 ;
        RECT 271.995 116.260 274.155 116.610 ;
        RECT 147.105 115.210 149.265 115.560 ;
        RECT 194.105 115.210 196.265 115.560 ;
        RECT 199.165 114.850 201.325 115.540 ;
        RECT 220.165 114.850 222.325 115.540 ;
        RECT 224.995 115.430 227.155 115.780 ;
        RECT 271.995 115.430 274.155 115.780 ;
        RECT 147.105 114.380 149.265 114.730 ;
        RECT 194.105 114.380 196.265 114.730 ;
        RECT 224.995 114.600 227.155 114.950 ;
        RECT 271.995 114.600 274.155 114.950 ;
        RECT 147.105 113.550 149.265 113.900 ;
        RECT 194.105 113.550 196.265 113.900 ;
        RECT 199.165 113.680 201.325 114.370 ;
        RECT 220.165 113.680 222.325 114.370 ;
        RECT 224.995 113.770 227.155 114.120 ;
        RECT 271.995 113.770 274.155 114.120 ;
        RECT 147.105 112.720 149.265 113.070 ;
        RECT 194.105 112.720 196.265 113.070 ;
        RECT 199.165 112.510 201.325 113.200 ;
        RECT 220.165 112.510 222.325 113.200 ;
        RECT 224.995 112.940 227.155 113.290 ;
        RECT 271.995 112.940 274.155 113.290 ;
        RECT 147.105 111.890 149.265 112.240 ;
        RECT 194.105 111.890 196.265 112.240 ;
        RECT 224.995 112.110 227.155 112.460 ;
        RECT 271.995 112.110 274.155 112.460 ;
        RECT 147.105 111.060 149.265 111.410 ;
        RECT 194.105 111.060 196.265 111.410 ;
        RECT 199.165 111.340 201.325 112.030 ;
        RECT 220.165 111.340 222.325 112.030 ;
        RECT 224.995 111.280 227.155 111.630 ;
        RECT 271.995 111.280 274.155 111.630 ;
        RECT 147.105 110.230 149.265 110.580 ;
        RECT 194.105 110.230 196.265 110.580 ;
        RECT 199.165 110.170 201.325 110.860 ;
        RECT 220.165 110.170 222.325 110.860 ;
        RECT 224.995 110.450 227.155 110.800 ;
        RECT 271.995 110.450 274.155 110.800 ;
        RECT 147.105 109.400 149.265 109.750 ;
        RECT 194.105 109.400 196.265 109.750 ;
        RECT 199.165 109.000 201.325 109.690 ;
        RECT 220.165 109.000 222.325 109.690 ;
        RECT 224.995 109.620 227.155 109.970 ;
        RECT 271.995 109.620 274.155 109.970 ;
        RECT 147.105 108.570 149.265 108.920 ;
        RECT 194.105 108.570 196.265 108.920 ;
        RECT 224.995 108.790 227.155 109.140 ;
        RECT 271.995 108.790 274.155 109.140 ;
        RECT 147.105 107.740 149.265 108.090 ;
        RECT 194.105 107.740 196.265 108.090 ;
        RECT 199.165 107.830 201.325 108.520 ;
        RECT 220.165 107.830 222.325 108.520 ;
        RECT 224.995 107.960 227.155 108.310 ;
        RECT 271.995 107.960 274.155 108.310 ;
        RECT 147.105 106.910 149.265 107.260 ;
        RECT 194.105 106.910 196.265 107.260 ;
        RECT 199.165 106.660 201.325 107.350 ;
        RECT 220.165 106.660 222.325 107.350 ;
        RECT 224.995 107.130 227.155 107.480 ;
        RECT 271.995 107.130 274.155 107.480 ;
        RECT 147.105 106.080 149.265 106.430 ;
        RECT 194.105 106.080 196.265 106.430 ;
        RECT 224.995 106.300 227.155 106.650 ;
        RECT 271.995 106.300 274.155 106.650 ;
        RECT 147.105 105.250 149.265 105.600 ;
        RECT 194.105 105.250 196.265 105.600 ;
        RECT 199.165 105.490 201.325 106.180 ;
        RECT 220.165 105.490 222.325 106.180 ;
        RECT 224.995 105.470 227.155 105.820 ;
        RECT 271.995 105.470 274.155 105.820 ;
        RECT 147.105 104.420 149.265 104.770 ;
        RECT 194.105 104.420 196.265 104.770 ;
        RECT 199.165 104.320 201.325 105.010 ;
        RECT 220.165 104.320 222.325 105.010 ;
        RECT 224.995 104.640 227.155 104.990 ;
        RECT 271.995 104.640 274.155 104.990 ;
        RECT 147.105 103.590 149.265 103.940 ;
        RECT 194.105 103.590 196.265 103.940 ;
        RECT 199.165 103.150 201.325 103.840 ;
        RECT 220.165 103.150 222.325 103.840 ;
        RECT 224.995 103.810 227.155 104.160 ;
        RECT 271.995 103.810 274.155 104.160 ;
        RECT 147.105 102.760 149.265 103.110 ;
        RECT 194.105 102.760 196.265 103.110 ;
        RECT 224.995 102.980 227.155 103.330 ;
        RECT 271.995 102.980 274.155 103.330 ;
        RECT 147.105 101.930 149.265 102.280 ;
        RECT 194.105 101.930 196.265 102.280 ;
        RECT 224.995 102.150 227.155 102.500 ;
        RECT 271.995 102.150 274.155 102.500 ;
        RECT 147.105 101.100 149.265 101.450 ;
        RECT 194.105 101.100 196.265 101.450 ;
        RECT 224.995 101.320 227.155 101.670 ;
        RECT 271.995 101.320 274.155 101.670 ;
        RECT 147.105 100.270 149.265 100.620 ;
        RECT 194.105 100.270 196.265 100.620 ;
        RECT 224.995 100.490 227.155 100.840 ;
        RECT 271.995 100.490 274.155 100.840 ;
        RECT 147.105 99.440 149.265 99.790 ;
        RECT 194.105 99.440 196.265 99.790 ;
        RECT 224.995 99.660 227.155 100.010 ;
        RECT 271.995 99.660 274.155 100.010 ;
        RECT 212.225 99.180 212.685 99.350 ;
        RECT 214.915 99.180 215.375 99.350 ;
        RECT 147.105 98.610 149.265 98.960 ;
        RECT 194.105 98.610 196.265 98.960 ;
        RECT 207.935 98.700 208.395 98.870 ;
        RECT 208.610 98.140 208.780 98.640 ;
        RECT 211.885 98.620 212.055 99.120 ;
        RECT 215.545 98.620 215.715 99.120 ;
        RECT 224.995 98.830 227.155 99.180 ;
        RECT 271.995 98.830 274.155 99.180 ;
        RECT 212.225 98.390 212.685 98.560 ;
        RECT 147.105 97.780 149.265 98.130 ;
        RECT 194.105 97.780 196.265 98.130 ;
        RECT 224.995 98.000 227.155 98.350 ;
        RECT 271.995 98.000 274.155 98.350 ;
        RECT 147.105 96.950 149.265 97.300 ;
        RECT 194.105 96.950 196.265 97.300 ;
        RECT 224.995 97.170 227.155 97.520 ;
        RECT 271.995 97.170 274.155 97.520 ;
        RECT 147.105 96.120 149.265 96.470 ;
        RECT 194.105 96.120 196.265 96.470 ;
        RECT 212.225 96.400 212.685 96.570 ;
        RECT 214.915 96.400 215.375 96.570 ;
        RECT 224.995 96.340 227.155 96.690 ;
        RECT 271.995 96.340 274.155 96.690 ;
        RECT 211.885 95.840 212.055 96.340 ;
        RECT 215.545 95.840 215.715 96.340 ;
        RECT 147.105 95.290 149.265 95.640 ;
        RECT 194.105 95.290 196.265 95.640 ;
        RECT 207.935 95.620 208.395 95.790 ;
        RECT 212.225 95.610 212.685 95.780 ;
        RECT 204.520 95.060 204.690 95.560 ;
        RECT 208.610 95.060 208.780 95.560 ;
        RECT 224.995 95.510 227.155 95.860 ;
        RECT 271.995 95.510 274.155 95.860 ;
        RECT 204.905 94.830 205.365 95.000 ;
        RECT 207.935 94.830 208.395 95.000 ;
        RECT 147.105 94.460 149.265 94.810 ;
        RECT 194.105 94.460 196.265 94.810 ;
        RECT 224.995 94.680 227.155 95.030 ;
        RECT 271.995 94.680 274.155 95.030 ;
        RECT 147.105 93.630 149.265 93.980 ;
        RECT 194.105 93.630 196.265 93.980 ;
        RECT 224.995 93.850 227.155 94.200 ;
        RECT 271.995 93.850 274.155 94.200 ;
        RECT 212.225 93.620 212.685 93.790 ;
        RECT 214.915 93.620 215.375 93.790 ;
        RECT 218.545 93.610 219.005 93.780 ;
        RECT 147.105 92.800 149.265 93.150 ;
        RECT 194.105 92.800 196.265 93.150 ;
        RECT 211.885 93.060 212.055 93.560 ;
        RECT 215.545 93.060 215.715 93.560 ;
        RECT 219.175 93.050 219.345 93.550 ;
        RECT 224.995 93.020 227.155 93.370 ;
        RECT 271.995 93.020 274.155 93.370 ;
        RECT 212.225 92.830 212.685 93.000 ;
        RECT 207.935 92.540 208.395 92.710 ;
        RECT 147.105 91.970 149.265 92.320 ;
        RECT 194.105 91.970 196.265 92.320 ;
        RECT 204.520 91.980 204.690 92.480 ;
        RECT 208.610 91.980 208.780 92.480 ;
        RECT 224.995 92.190 227.155 92.540 ;
        RECT 271.995 92.190 274.155 92.540 ;
        RECT 204.905 91.750 205.365 91.920 ;
        RECT 207.935 91.750 208.395 91.920 ;
        RECT 147.105 91.140 149.265 91.490 ;
        RECT 194.105 91.140 196.265 91.490 ;
        RECT 224.995 91.360 227.155 91.710 ;
        RECT 271.995 91.360 274.155 91.710 ;
        RECT 212.225 90.840 212.685 91.010 ;
        RECT 214.915 90.840 215.375 91.010 ;
        RECT 147.105 90.310 149.265 90.660 ;
        RECT 194.105 90.310 196.265 90.660 ;
        RECT 215.545 90.280 215.715 90.780 ;
        RECT 219.175 90.270 219.345 90.770 ;
        RECT 224.995 90.530 227.155 90.880 ;
        RECT 271.995 90.530 274.155 90.880 ;
        RECT 212.225 90.050 212.685 90.220 ;
        RECT 147.105 89.480 149.265 89.830 ;
        RECT 194.105 89.480 196.265 89.830 ;
        RECT 224.995 89.700 227.155 90.050 ;
        RECT 271.995 89.700 274.155 90.050 ;
        RECT 207.935 89.460 208.395 89.630 ;
        RECT 147.105 88.650 149.265 89.000 ;
        RECT 194.105 88.650 196.265 89.000 ;
        RECT 204.520 88.900 204.690 89.400 ;
        RECT 224.995 88.870 227.155 89.220 ;
        RECT 271.995 88.870 274.155 89.220 ;
        RECT 204.905 88.670 205.365 88.840 ;
        RECT 207.935 88.670 208.395 88.840 ;
        RECT 147.105 87.820 149.265 88.170 ;
        RECT 194.105 87.820 196.265 88.170 ;
        RECT 212.225 88.060 212.685 88.230 ;
        RECT 214.915 88.060 215.375 88.230 ;
        RECT 218.545 88.050 219.005 88.220 ;
        RECT 224.995 88.040 227.155 88.390 ;
        RECT 271.995 88.040 274.155 88.390 ;
        RECT 211.885 87.500 212.055 88.000 ;
        RECT 215.545 87.500 215.715 88.000 ;
        RECT 219.175 87.490 219.345 87.990 ;
        RECT 147.105 86.990 149.265 87.340 ;
        RECT 194.105 86.990 196.265 87.340 ;
        RECT 212.225 87.270 212.685 87.440 ;
        RECT 224.995 87.210 227.155 87.560 ;
        RECT 271.995 87.210 274.155 87.560 ;
        RECT 147.105 86.160 149.265 86.510 ;
        RECT 194.105 86.160 196.265 86.510 ;
        RECT 204.905 86.380 205.365 86.550 ;
        RECT 207.935 86.380 208.395 86.550 ;
        RECT 224.995 86.380 227.155 86.730 ;
        RECT 271.995 86.380 274.155 86.730 ;
        RECT 204.520 85.820 204.690 86.320 ;
        RECT 208.610 85.820 208.780 86.320 ;
        RECT 147.105 85.330 149.265 85.680 ;
        RECT 194.105 85.330 196.265 85.680 ;
        RECT 224.995 85.550 227.155 85.900 ;
        RECT 271.995 85.550 274.155 85.900 ;
        RECT 212.225 85.280 212.685 85.450 ;
        RECT 214.915 85.280 215.375 85.450 ;
        RECT 218.545 85.270 219.005 85.440 ;
        RECT 194.105 84.500 196.265 84.850 ;
        RECT 211.885 84.720 212.055 85.220 ;
        RECT 215.545 84.720 215.715 85.220 ;
        RECT 219.175 84.710 219.345 85.210 ;
        RECT 224.995 84.720 227.155 85.070 ;
        RECT 271.995 84.720 274.155 85.070 ;
        RECT 212.225 84.490 212.685 84.660 ;
        RECT 218.545 84.480 219.005 84.650 ;
        RECT 224.995 83.890 227.155 84.240 ;
        RECT 271.995 83.890 274.155 84.240 ;
        RECT 224.995 83.060 227.155 83.410 ;
        RECT 271.995 83.060 274.155 83.410 ;
        RECT 224.995 82.230 227.155 82.580 ;
        RECT 271.995 82.230 274.155 82.580 ;
        RECT 147.155 81.500 149.315 81.850 ;
        RECT 194.155 81.500 196.315 81.850 ;
        RECT 224.995 81.400 227.155 81.750 ;
        RECT 271.995 81.400 274.155 81.750 ;
        RECT 147.155 80.670 149.315 81.020 ;
        RECT 194.155 80.670 196.315 81.020 ;
        RECT 224.995 80.570 227.155 80.920 ;
        RECT 271.995 80.570 274.155 80.920 ;
        RECT 147.155 79.840 149.315 80.190 ;
        RECT 194.155 79.840 196.315 80.190 ;
        RECT 147.155 79.010 149.315 79.360 ;
        RECT 194.155 79.010 196.315 79.360 ;
        RECT 147.155 78.180 149.315 78.530 ;
        RECT 194.155 78.180 196.315 78.530 ;
        RECT 147.155 77.350 149.315 77.700 ;
        RECT 194.155 77.350 196.315 77.700 ;
        RECT 147.155 76.520 149.315 76.870 ;
        RECT 194.155 76.520 196.315 76.870 ;
        RECT 147.155 75.690 149.315 76.040 ;
        RECT 194.155 75.690 196.315 76.040 ;
        RECT 147.155 74.860 149.315 75.210 ;
        RECT 194.155 74.860 196.315 75.210 ;
        RECT 198.910 74.600 199.390 80.290 ;
        RECT 204.955 79.100 205.415 79.270 ;
        RECT 208.305 79.100 208.765 79.270 ;
        RECT 212.815 79.100 213.275 79.270 ;
        RECT 216.165 79.100 216.625 79.270 ;
        RECT 201.120 78.530 201.290 79.030 ;
        RECT 202.090 78.530 202.260 79.030 ;
        RECT 204.570 78.540 204.740 79.040 ;
        RECT 205.630 78.540 205.800 79.040 ;
        RECT 207.920 78.540 208.090 79.040 ;
        RECT 208.980 78.540 209.150 79.040 ;
        RECT 212.430 78.540 212.600 79.040 ;
        RECT 213.490 78.540 213.660 79.040 ;
        RECT 215.780 78.540 215.950 79.040 ;
        RECT 216.840 78.540 217.010 79.040 ;
        RECT 219.320 78.530 219.490 79.030 ;
        RECT 220.290 78.530 220.460 79.030 ;
        RECT 201.460 78.300 201.920 78.470 ;
        RECT 204.955 78.310 205.415 78.480 ;
        RECT 216.165 78.310 216.625 78.480 ;
        RECT 219.660 78.300 220.120 78.470 ;
        RECT 201.450 76.060 201.910 76.230 ;
        RECT 204.965 76.050 205.425 76.220 ;
        RECT 216.155 76.050 216.615 76.220 ;
        RECT 219.670 76.060 220.130 76.230 ;
        RECT 204.580 75.490 204.750 75.990 ;
        RECT 205.640 75.490 205.810 75.990 ;
        RECT 207.920 75.460 208.090 75.960 ;
        RECT 208.980 75.460 209.150 75.960 ;
        RECT 212.430 75.460 212.600 75.960 ;
        RECT 213.490 75.460 213.660 75.960 ;
        RECT 215.770 75.490 215.940 75.990 ;
        RECT 216.830 75.490 217.000 75.990 ;
        RECT 204.965 75.260 205.425 75.430 ;
        RECT 208.305 75.230 208.765 75.400 ;
        RECT 212.815 75.230 213.275 75.400 ;
        RECT 216.155 75.260 216.615 75.430 ;
        RECT 222.190 74.600 222.670 80.290 ;
        RECT 224.995 79.740 227.155 80.090 ;
        RECT 271.995 79.740 274.155 80.090 ;
        RECT 224.995 78.910 227.155 79.260 ;
        RECT 271.995 78.910 274.155 79.260 ;
        RECT 224.995 78.080 227.155 78.430 ;
        RECT 271.995 78.080 274.155 78.430 ;
        RECT 224.995 77.250 227.155 77.600 ;
        RECT 271.995 77.250 274.155 77.600 ;
        RECT 224.995 76.420 227.155 76.770 ;
        RECT 271.995 76.420 274.155 76.770 ;
        RECT 224.995 75.590 227.155 75.940 ;
        RECT 271.995 75.590 274.155 75.940 ;
        RECT 224.995 74.760 227.155 75.110 ;
        RECT 271.995 74.760 274.155 75.110 ;
        RECT 147.155 74.030 149.315 74.380 ;
        RECT 194.155 74.030 196.315 74.380 ;
        RECT 224.995 73.930 227.155 74.280 ;
        RECT 271.995 73.930 274.155 74.280 ;
        RECT 147.155 73.200 149.315 73.550 ;
        RECT 194.155 73.200 196.315 73.550 ;
        RECT 224.995 73.100 227.155 73.450 ;
        RECT 271.995 73.100 274.155 73.450 ;
        RECT 147.155 72.370 149.315 72.720 ;
        RECT 194.155 72.370 196.315 72.720 ;
        RECT 224.995 72.270 227.155 72.620 ;
        RECT 271.995 72.270 274.155 72.620 ;
        RECT 147.155 71.540 149.315 71.890 ;
        RECT 194.155 71.540 196.315 71.890 ;
        RECT 224.995 71.440 227.155 71.790 ;
        RECT 271.995 71.440 274.155 71.790 ;
        RECT 147.155 70.710 149.315 71.060 ;
        RECT 194.155 70.710 196.315 71.060 ;
        RECT 215.795 70.320 217.955 71.010 ;
        RECT 224.995 70.610 227.155 70.960 ;
        RECT 271.995 70.610 274.155 70.960 ;
        RECT 147.155 69.880 149.315 70.230 ;
        RECT 194.155 69.880 196.315 70.230 ;
        RECT 224.995 69.780 227.155 70.130 ;
        RECT 271.995 69.780 274.155 70.130 ;
        RECT 147.155 69.050 149.315 69.400 ;
        RECT 194.155 69.050 196.315 69.400 ;
        RECT 224.995 68.950 227.155 69.300 ;
        RECT 271.995 68.950 274.155 69.300 ;
        RECT 147.155 68.220 149.315 68.570 ;
        RECT 194.155 68.220 196.315 68.570 ;
        RECT 224.995 68.120 227.155 68.470 ;
        RECT 271.995 68.120 274.155 68.470 ;
        RECT 147.155 67.390 149.315 67.740 ;
        RECT 194.155 67.390 196.315 67.740 ;
        RECT 202.780 67.610 203.820 67.780 ;
        RECT 205.970 67.610 207.010 67.780 ;
        RECT 214.570 67.610 215.610 67.780 ;
        RECT 217.760 67.610 218.800 67.780 ;
        RECT 224.995 67.290 227.155 67.640 ;
        RECT 271.995 67.290 274.155 67.640 ;
        RECT 194.155 66.560 196.315 66.910 ;
        RECT 209.655 66.885 209.825 67.215 ;
        RECT 209.995 66.745 210.535 66.915 ;
        RECT 224.995 66.460 227.155 66.810 ;
        RECT 271.995 66.460 274.155 66.810 ;
        RECT 205.655 64.680 206.695 64.850 ;
        RECT 206.910 64.820 207.080 65.150 ;
        RECT 209.995 65.120 210.535 65.290 ;
        RECT 209.995 64.680 210.535 64.850 ;
        RECT 211.945 64.820 212.115 65.150 ;
        RECT 212.285 64.680 212.745 64.850 ;
      LAYER mcon ;
        RECT 147.205 131.070 147.375 131.240 ;
        RECT 147.565 131.070 147.735 131.240 ;
        RECT 147.925 131.070 148.095 131.240 ;
        RECT 148.285 131.070 148.455 131.240 ;
        RECT 148.645 131.070 148.815 131.240 ;
        RECT 149.005 131.070 149.175 131.240 ;
        RECT 194.200 131.070 194.370 131.240 ;
        RECT 194.560 131.070 194.730 131.240 ;
        RECT 194.920 131.070 195.090 131.240 ;
        RECT 195.280 131.070 195.450 131.240 ;
        RECT 195.640 131.070 195.810 131.240 ;
        RECT 196.000 131.070 196.170 131.240 ;
        RECT 225.095 131.290 225.265 131.460 ;
        RECT 225.455 131.290 225.625 131.460 ;
        RECT 225.815 131.290 225.985 131.460 ;
        RECT 226.175 131.290 226.345 131.460 ;
        RECT 226.535 131.290 226.705 131.460 ;
        RECT 226.895 131.290 227.065 131.460 ;
        RECT 147.205 130.240 147.375 130.410 ;
        RECT 147.565 130.240 147.735 130.410 ;
        RECT 147.925 130.240 148.095 130.410 ;
        RECT 148.285 130.240 148.455 130.410 ;
        RECT 148.645 130.240 148.815 130.410 ;
        RECT 149.005 130.240 149.175 130.410 ;
        RECT 194.200 130.240 194.370 130.410 ;
        RECT 194.560 130.240 194.730 130.410 ;
        RECT 194.920 130.240 195.090 130.410 ;
        RECT 195.280 130.240 195.450 130.410 ;
        RECT 195.640 130.240 195.810 130.410 ;
        RECT 196.000 130.240 196.170 130.410 ;
        RECT 199.265 130.140 201.235 130.670 ;
        RECT 225.095 130.460 225.265 130.630 ;
        RECT 225.455 130.460 225.625 130.630 ;
        RECT 225.815 130.460 225.985 130.630 ;
        RECT 226.175 130.460 226.345 130.630 ;
        RECT 226.535 130.460 226.705 130.630 ;
        RECT 226.895 130.460 227.065 130.630 ;
        RECT 272.090 130.460 272.260 130.630 ;
        RECT 272.450 130.460 272.620 130.630 ;
        RECT 272.810 130.460 272.980 130.630 ;
        RECT 273.170 130.460 273.340 130.630 ;
        RECT 273.530 130.460 273.700 130.630 ;
        RECT 273.890 130.460 274.060 130.630 ;
        RECT 147.205 129.410 147.375 129.580 ;
        RECT 147.565 129.410 147.735 129.580 ;
        RECT 147.925 129.410 148.095 129.580 ;
        RECT 148.285 129.410 148.455 129.580 ;
        RECT 148.645 129.410 148.815 129.580 ;
        RECT 149.005 129.410 149.175 129.580 ;
        RECT 225.095 129.630 225.265 129.800 ;
        RECT 225.455 129.630 225.625 129.800 ;
        RECT 225.815 129.630 225.985 129.800 ;
        RECT 226.175 129.630 226.345 129.800 ;
        RECT 226.535 129.630 226.705 129.800 ;
        RECT 226.895 129.630 227.065 129.800 ;
        RECT 194.200 129.410 194.370 129.580 ;
        RECT 194.560 129.410 194.730 129.580 ;
        RECT 194.920 129.410 195.090 129.580 ;
        RECT 195.280 129.410 195.450 129.580 ;
        RECT 195.640 129.410 195.810 129.580 ;
        RECT 196.000 129.410 196.170 129.580 ;
        RECT 199.265 128.970 201.235 129.500 ;
        RECT 272.090 129.630 272.260 129.800 ;
        RECT 272.450 129.630 272.620 129.800 ;
        RECT 272.810 129.630 272.980 129.800 ;
        RECT 273.170 129.630 273.340 129.800 ;
        RECT 273.530 129.630 273.700 129.800 ;
        RECT 273.890 129.630 274.060 129.800 ;
        RECT 220.260 128.970 222.230 129.500 ;
        RECT 147.205 128.580 147.375 128.750 ;
        RECT 147.565 128.580 147.735 128.750 ;
        RECT 147.925 128.580 148.095 128.750 ;
        RECT 148.285 128.580 148.455 128.750 ;
        RECT 148.645 128.580 148.815 128.750 ;
        RECT 149.005 128.580 149.175 128.750 ;
        RECT 194.200 128.580 194.370 128.750 ;
        RECT 194.560 128.580 194.730 128.750 ;
        RECT 194.920 128.580 195.090 128.750 ;
        RECT 195.280 128.580 195.450 128.750 ;
        RECT 195.640 128.580 195.810 128.750 ;
        RECT 196.000 128.580 196.170 128.750 ;
        RECT 225.095 128.800 225.265 128.970 ;
        RECT 225.455 128.800 225.625 128.970 ;
        RECT 225.815 128.800 225.985 128.970 ;
        RECT 226.175 128.800 226.345 128.970 ;
        RECT 226.535 128.800 226.705 128.970 ;
        RECT 226.895 128.800 227.065 128.970 ;
        RECT 272.090 128.800 272.260 128.970 ;
        RECT 272.450 128.800 272.620 128.970 ;
        RECT 272.810 128.800 272.980 128.970 ;
        RECT 273.170 128.800 273.340 128.970 ;
        RECT 273.530 128.800 273.700 128.970 ;
        RECT 273.890 128.800 274.060 128.970 ;
        RECT 147.205 127.750 147.375 127.920 ;
        RECT 147.565 127.750 147.735 127.920 ;
        RECT 147.925 127.750 148.095 127.920 ;
        RECT 148.285 127.750 148.455 127.920 ;
        RECT 148.645 127.750 148.815 127.920 ;
        RECT 149.005 127.750 149.175 127.920 ;
        RECT 194.200 127.750 194.370 127.920 ;
        RECT 194.560 127.750 194.730 127.920 ;
        RECT 194.920 127.750 195.090 127.920 ;
        RECT 195.280 127.750 195.450 127.920 ;
        RECT 195.640 127.750 195.810 127.920 ;
        RECT 196.000 127.750 196.170 127.920 ;
        RECT 199.265 127.800 201.235 128.330 ;
        RECT 220.260 127.800 222.230 128.330 ;
        RECT 225.095 127.970 225.265 128.140 ;
        RECT 225.455 127.970 225.625 128.140 ;
        RECT 225.815 127.970 225.985 128.140 ;
        RECT 226.175 127.970 226.345 128.140 ;
        RECT 226.535 127.970 226.705 128.140 ;
        RECT 226.895 127.970 227.065 128.140 ;
        RECT 272.090 127.970 272.260 128.140 ;
        RECT 272.450 127.970 272.620 128.140 ;
        RECT 272.810 127.970 272.980 128.140 ;
        RECT 273.170 127.970 273.340 128.140 ;
        RECT 273.530 127.970 273.700 128.140 ;
        RECT 273.890 127.970 274.060 128.140 ;
        RECT 147.205 126.920 147.375 127.090 ;
        RECT 147.565 126.920 147.735 127.090 ;
        RECT 147.925 126.920 148.095 127.090 ;
        RECT 148.285 126.920 148.455 127.090 ;
        RECT 148.645 126.920 148.815 127.090 ;
        RECT 149.005 126.920 149.175 127.090 ;
        RECT 194.200 126.920 194.370 127.090 ;
        RECT 194.560 126.920 194.730 127.090 ;
        RECT 194.920 126.920 195.090 127.090 ;
        RECT 195.280 126.920 195.450 127.090 ;
        RECT 195.640 126.920 195.810 127.090 ;
        RECT 196.000 126.920 196.170 127.090 ;
        RECT 199.265 126.630 201.235 127.160 ;
        RECT 220.260 126.630 222.230 127.160 ;
        RECT 225.095 127.140 225.265 127.310 ;
        RECT 225.455 127.140 225.625 127.310 ;
        RECT 225.815 127.140 225.985 127.310 ;
        RECT 226.175 127.140 226.345 127.310 ;
        RECT 226.535 127.140 226.705 127.310 ;
        RECT 226.895 127.140 227.065 127.310 ;
        RECT 272.090 127.140 272.260 127.310 ;
        RECT 272.450 127.140 272.620 127.310 ;
        RECT 272.810 127.140 272.980 127.310 ;
        RECT 273.170 127.140 273.340 127.310 ;
        RECT 273.530 127.140 273.700 127.310 ;
        RECT 273.890 127.140 274.060 127.310 ;
        RECT 147.205 126.090 147.375 126.260 ;
        RECT 147.565 126.090 147.735 126.260 ;
        RECT 147.925 126.090 148.095 126.260 ;
        RECT 148.285 126.090 148.455 126.260 ;
        RECT 148.645 126.090 148.815 126.260 ;
        RECT 149.005 126.090 149.175 126.260 ;
        RECT 194.200 126.090 194.370 126.260 ;
        RECT 194.560 126.090 194.730 126.260 ;
        RECT 194.920 126.090 195.090 126.260 ;
        RECT 195.280 126.090 195.450 126.260 ;
        RECT 195.640 126.090 195.810 126.260 ;
        RECT 196.000 126.090 196.170 126.260 ;
        RECT 225.095 126.310 225.265 126.480 ;
        RECT 225.455 126.310 225.625 126.480 ;
        RECT 225.815 126.310 225.985 126.480 ;
        RECT 226.175 126.310 226.345 126.480 ;
        RECT 226.535 126.310 226.705 126.480 ;
        RECT 226.895 126.310 227.065 126.480 ;
        RECT 272.090 126.310 272.260 126.480 ;
        RECT 272.450 126.310 272.620 126.480 ;
        RECT 272.810 126.310 272.980 126.480 ;
        RECT 273.170 126.310 273.340 126.480 ;
        RECT 273.530 126.310 273.700 126.480 ;
        RECT 273.890 126.310 274.060 126.480 ;
        RECT 147.205 125.260 147.375 125.430 ;
        RECT 147.565 125.260 147.735 125.430 ;
        RECT 147.925 125.260 148.095 125.430 ;
        RECT 148.285 125.260 148.455 125.430 ;
        RECT 148.645 125.260 148.815 125.430 ;
        RECT 149.005 125.260 149.175 125.430 ;
        RECT 194.200 125.260 194.370 125.430 ;
        RECT 194.560 125.260 194.730 125.430 ;
        RECT 194.920 125.260 195.090 125.430 ;
        RECT 195.280 125.260 195.450 125.430 ;
        RECT 195.640 125.260 195.810 125.430 ;
        RECT 196.000 125.260 196.170 125.430 ;
        RECT 199.265 125.460 201.235 125.990 ;
        RECT 220.260 125.460 222.230 125.990 ;
        RECT 225.095 125.480 225.265 125.650 ;
        RECT 225.455 125.480 225.625 125.650 ;
        RECT 225.815 125.480 225.985 125.650 ;
        RECT 226.175 125.480 226.345 125.650 ;
        RECT 226.535 125.480 226.705 125.650 ;
        RECT 226.895 125.480 227.065 125.650 ;
        RECT 272.090 125.480 272.260 125.650 ;
        RECT 272.450 125.480 272.620 125.650 ;
        RECT 272.810 125.480 272.980 125.650 ;
        RECT 273.170 125.480 273.340 125.650 ;
        RECT 273.530 125.480 273.700 125.650 ;
        RECT 273.890 125.480 274.060 125.650 ;
        RECT 147.205 124.430 147.375 124.600 ;
        RECT 147.565 124.430 147.735 124.600 ;
        RECT 147.925 124.430 148.095 124.600 ;
        RECT 148.285 124.430 148.455 124.600 ;
        RECT 148.645 124.430 148.815 124.600 ;
        RECT 149.005 124.430 149.175 124.600 ;
        RECT 194.200 124.430 194.370 124.600 ;
        RECT 194.560 124.430 194.730 124.600 ;
        RECT 194.920 124.430 195.090 124.600 ;
        RECT 195.280 124.430 195.450 124.600 ;
        RECT 195.640 124.430 195.810 124.600 ;
        RECT 196.000 124.430 196.170 124.600 ;
        RECT 199.265 124.290 201.235 124.820 ;
        RECT 220.260 124.290 222.230 124.820 ;
        RECT 225.095 124.650 225.265 124.820 ;
        RECT 225.455 124.650 225.625 124.820 ;
        RECT 225.815 124.650 225.985 124.820 ;
        RECT 226.175 124.650 226.345 124.820 ;
        RECT 226.535 124.650 226.705 124.820 ;
        RECT 226.895 124.650 227.065 124.820 ;
        RECT 272.090 124.650 272.260 124.820 ;
        RECT 272.450 124.650 272.620 124.820 ;
        RECT 272.810 124.650 272.980 124.820 ;
        RECT 273.170 124.650 273.340 124.820 ;
        RECT 273.530 124.650 273.700 124.820 ;
        RECT 273.890 124.650 274.060 124.820 ;
        RECT 147.205 123.600 147.375 123.770 ;
        RECT 147.565 123.600 147.735 123.770 ;
        RECT 147.925 123.600 148.095 123.770 ;
        RECT 148.285 123.600 148.455 123.770 ;
        RECT 148.645 123.600 148.815 123.770 ;
        RECT 149.005 123.600 149.175 123.770 ;
        RECT 194.200 123.600 194.370 123.770 ;
        RECT 194.560 123.600 194.730 123.770 ;
        RECT 194.920 123.600 195.090 123.770 ;
        RECT 195.280 123.600 195.450 123.770 ;
        RECT 195.640 123.600 195.810 123.770 ;
        RECT 196.000 123.600 196.170 123.770 ;
        RECT 225.095 123.820 225.265 123.990 ;
        RECT 225.455 123.820 225.625 123.990 ;
        RECT 225.815 123.820 225.985 123.990 ;
        RECT 226.175 123.820 226.345 123.990 ;
        RECT 226.535 123.820 226.705 123.990 ;
        RECT 226.895 123.820 227.065 123.990 ;
        RECT 272.090 123.820 272.260 123.990 ;
        RECT 272.450 123.820 272.620 123.990 ;
        RECT 272.810 123.820 272.980 123.990 ;
        RECT 273.170 123.820 273.340 123.990 ;
        RECT 273.530 123.820 273.700 123.990 ;
        RECT 273.890 123.820 274.060 123.990 ;
        RECT 199.265 123.120 201.235 123.650 ;
        RECT 220.260 123.120 222.230 123.650 ;
        RECT 147.205 122.770 147.375 122.940 ;
        RECT 147.565 122.770 147.735 122.940 ;
        RECT 147.925 122.770 148.095 122.940 ;
        RECT 148.285 122.770 148.455 122.940 ;
        RECT 148.645 122.770 148.815 122.940 ;
        RECT 149.005 122.770 149.175 122.940 ;
        RECT 194.200 122.770 194.370 122.940 ;
        RECT 194.560 122.770 194.730 122.940 ;
        RECT 194.920 122.770 195.090 122.940 ;
        RECT 195.280 122.770 195.450 122.940 ;
        RECT 195.640 122.770 195.810 122.940 ;
        RECT 196.000 122.770 196.170 122.940 ;
        RECT 225.095 122.990 225.265 123.160 ;
        RECT 225.455 122.990 225.625 123.160 ;
        RECT 225.815 122.990 225.985 123.160 ;
        RECT 226.175 122.990 226.345 123.160 ;
        RECT 226.535 122.990 226.705 123.160 ;
        RECT 226.895 122.990 227.065 123.160 ;
        RECT 272.090 122.990 272.260 123.160 ;
        RECT 272.450 122.990 272.620 123.160 ;
        RECT 272.810 122.990 272.980 123.160 ;
        RECT 273.170 122.990 273.340 123.160 ;
        RECT 273.530 122.990 273.700 123.160 ;
        RECT 273.890 122.990 274.060 123.160 ;
        RECT 147.205 121.940 147.375 122.110 ;
        RECT 147.565 121.940 147.735 122.110 ;
        RECT 147.925 121.940 148.095 122.110 ;
        RECT 148.285 121.940 148.455 122.110 ;
        RECT 148.645 121.940 148.815 122.110 ;
        RECT 149.005 121.940 149.175 122.110 ;
        RECT 194.200 121.940 194.370 122.110 ;
        RECT 194.560 121.940 194.730 122.110 ;
        RECT 194.920 121.940 195.090 122.110 ;
        RECT 195.280 121.940 195.450 122.110 ;
        RECT 195.640 121.940 195.810 122.110 ;
        RECT 196.000 121.940 196.170 122.110 ;
        RECT 199.265 121.950 201.235 122.480 ;
        RECT 220.260 121.950 222.230 122.480 ;
        RECT 225.095 122.160 225.265 122.330 ;
        RECT 225.455 122.160 225.625 122.330 ;
        RECT 225.815 122.160 225.985 122.330 ;
        RECT 226.175 122.160 226.345 122.330 ;
        RECT 226.535 122.160 226.705 122.330 ;
        RECT 226.895 122.160 227.065 122.330 ;
        RECT 272.090 122.160 272.260 122.330 ;
        RECT 272.450 122.160 272.620 122.330 ;
        RECT 272.810 122.160 272.980 122.330 ;
        RECT 273.170 122.160 273.340 122.330 ;
        RECT 273.530 122.160 273.700 122.330 ;
        RECT 273.890 122.160 274.060 122.330 ;
        RECT 147.205 121.110 147.375 121.280 ;
        RECT 147.565 121.110 147.735 121.280 ;
        RECT 147.925 121.110 148.095 121.280 ;
        RECT 148.285 121.110 148.455 121.280 ;
        RECT 148.645 121.110 148.815 121.280 ;
        RECT 149.005 121.110 149.175 121.280 ;
        RECT 194.200 121.110 194.370 121.280 ;
        RECT 194.560 121.110 194.730 121.280 ;
        RECT 194.920 121.110 195.090 121.280 ;
        RECT 195.280 121.110 195.450 121.280 ;
        RECT 195.640 121.110 195.810 121.280 ;
        RECT 196.000 121.110 196.170 121.280 ;
        RECT 199.265 120.780 201.235 121.310 ;
        RECT 220.260 120.780 222.230 121.310 ;
        RECT 225.095 121.330 225.265 121.500 ;
        RECT 225.455 121.330 225.625 121.500 ;
        RECT 225.815 121.330 225.985 121.500 ;
        RECT 226.175 121.330 226.345 121.500 ;
        RECT 226.535 121.330 226.705 121.500 ;
        RECT 226.895 121.330 227.065 121.500 ;
        RECT 272.090 121.330 272.260 121.500 ;
        RECT 272.450 121.330 272.620 121.500 ;
        RECT 272.810 121.330 272.980 121.500 ;
        RECT 273.170 121.330 273.340 121.500 ;
        RECT 273.530 121.330 273.700 121.500 ;
        RECT 273.890 121.330 274.060 121.500 ;
        RECT 147.205 120.280 147.375 120.450 ;
        RECT 147.565 120.280 147.735 120.450 ;
        RECT 147.925 120.280 148.095 120.450 ;
        RECT 148.285 120.280 148.455 120.450 ;
        RECT 148.645 120.280 148.815 120.450 ;
        RECT 149.005 120.280 149.175 120.450 ;
        RECT 194.200 120.280 194.370 120.450 ;
        RECT 194.560 120.280 194.730 120.450 ;
        RECT 194.920 120.280 195.090 120.450 ;
        RECT 195.280 120.280 195.450 120.450 ;
        RECT 195.640 120.280 195.810 120.450 ;
        RECT 196.000 120.280 196.170 120.450 ;
        RECT 225.095 120.500 225.265 120.670 ;
        RECT 225.455 120.500 225.625 120.670 ;
        RECT 225.815 120.500 225.985 120.670 ;
        RECT 226.175 120.500 226.345 120.670 ;
        RECT 226.535 120.500 226.705 120.670 ;
        RECT 226.895 120.500 227.065 120.670 ;
        RECT 272.090 120.500 272.260 120.670 ;
        RECT 272.450 120.500 272.620 120.670 ;
        RECT 272.810 120.500 272.980 120.670 ;
        RECT 273.170 120.500 273.340 120.670 ;
        RECT 273.530 120.500 273.700 120.670 ;
        RECT 273.890 120.500 274.060 120.670 ;
        RECT 147.205 119.450 147.375 119.620 ;
        RECT 147.565 119.450 147.735 119.620 ;
        RECT 147.925 119.450 148.095 119.620 ;
        RECT 148.285 119.450 148.455 119.620 ;
        RECT 148.645 119.450 148.815 119.620 ;
        RECT 149.005 119.450 149.175 119.620 ;
        RECT 194.200 119.450 194.370 119.620 ;
        RECT 194.560 119.450 194.730 119.620 ;
        RECT 194.920 119.450 195.090 119.620 ;
        RECT 195.280 119.450 195.450 119.620 ;
        RECT 195.640 119.450 195.810 119.620 ;
        RECT 196.000 119.450 196.170 119.620 ;
        RECT 199.265 119.610 201.235 120.140 ;
        RECT 220.260 119.610 222.230 120.140 ;
        RECT 225.095 119.670 225.265 119.840 ;
        RECT 225.455 119.670 225.625 119.840 ;
        RECT 225.815 119.670 225.985 119.840 ;
        RECT 226.175 119.670 226.345 119.840 ;
        RECT 226.535 119.670 226.705 119.840 ;
        RECT 226.895 119.670 227.065 119.840 ;
        RECT 272.090 119.670 272.260 119.840 ;
        RECT 272.450 119.670 272.620 119.840 ;
        RECT 272.810 119.670 272.980 119.840 ;
        RECT 273.170 119.670 273.340 119.840 ;
        RECT 273.530 119.670 273.700 119.840 ;
        RECT 273.890 119.670 274.060 119.840 ;
        RECT 147.205 118.620 147.375 118.790 ;
        RECT 147.565 118.620 147.735 118.790 ;
        RECT 147.925 118.620 148.095 118.790 ;
        RECT 148.285 118.620 148.455 118.790 ;
        RECT 148.645 118.620 148.815 118.790 ;
        RECT 149.005 118.620 149.175 118.790 ;
        RECT 194.200 118.620 194.370 118.790 ;
        RECT 194.560 118.620 194.730 118.790 ;
        RECT 194.920 118.620 195.090 118.790 ;
        RECT 195.280 118.620 195.450 118.790 ;
        RECT 195.640 118.620 195.810 118.790 ;
        RECT 196.000 118.620 196.170 118.790 ;
        RECT 199.265 118.440 201.235 118.970 ;
        RECT 220.260 118.440 222.230 118.970 ;
        RECT 225.095 118.840 225.265 119.010 ;
        RECT 225.455 118.840 225.625 119.010 ;
        RECT 225.815 118.840 225.985 119.010 ;
        RECT 226.175 118.840 226.345 119.010 ;
        RECT 226.535 118.840 226.705 119.010 ;
        RECT 226.895 118.840 227.065 119.010 ;
        RECT 272.090 118.840 272.260 119.010 ;
        RECT 272.450 118.840 272.620 119.010 ;
        RECT 272.810 118.840 272.980 119.010 ;
        RECT 273.170 118.840 273.340 119.010 ;
        RECT 273.530 118.840 273.700 119.010 ;
        RECT 273.890 118.840 274.060 119.010 ;
        RECT 147.205 117.790 147.375 117.960 ;
        RECT 147.565 117.790 147.735 117.960 ;
        RECT 147.925 117.790 148.095 117.960 ;
        RECT 148.285 117.790 148.455 117.960 ;
        RECT 148.645 117.790 148.815 117.960 ;
        RECT 149.005 117.790 149.175 117.960 ;
        RECT 194.200 117.790 194.370 117.960 ;
        RECT 194.560 117.790 194.730 117.960 ;
        RECT 194.920 117.790 195.090 117.960 ;
        RECT 195.280 117.790 195.450 117.960 ;
        RECT 195.640 117.790 195.810 117.960 ;
        RECT 196.000 117.790 196.170 117.960 ;
        RECT 225.095 118.010 225.265 118.180 ;
        RECT 225.455 118.010 225.625 118.180 ;
        RECT 225.815 118.010 225.985 118.180 ;
        RECT 226.175 118.010 226.345 118.180 ;
        RECT 226.535 118.010 226.705 118.180 ;
        RECT 226.895 118.010 227.065 118.180 ;
        RECT 272.090 118.010 272.260 118.180 ;
        RECT 272.450 118.010 272.620 118.180 ;
        RECT 272.810 118.010 272.980 118.180 ;
        RECT 273.170 118.010 273.340 118.180 ;
        RECT 273.530 118.010 273.700 118.180 ;
        RECT 273.890 118.010 274.060 118.180 ;
        RECT 199.265 117.270 201.235 117.800 ;
        RECT 147.205 116.960 147.375 117.130 ;
        RECT 147.565 116.960 147.735 117.130 ;
        RECT 147.925 116.960 148.095 117.130 ;
        RECT 148.285 116.960 148.455 117.130 ;
        RECT 148.645 116.960 148.815 117.130 ;
        RECT 149.005 116.960 149.175 117.130 ;
        RECT 220.260 117.270 222.230 117.800 ;
        RECT 194.200 116.960 194.370 117.130 ;
        RECT 194.560 116.960 194.730 117.130 ;
        RECT 194.920 116.960 195.090 117.130 ;
        RECT 195.280 116.960 195.450 117.130 ;
        RECT 195.640 116.960 195.810 117.130 ;
        RECT 196.000 116.960 196.170 117.130 ;
        RECT 225.095 117.180 225.265 117.350 ;
        RECT 225.455 117.180 225.625 117.350 ;
        RECT 225.815 117.180 225.985 117.350 ;
        RECT 226.175 117.180 226.345 117.350 ;
        RECT 226.535 117.180 226.705 117.350 ;
        RECT 226.895 117.180 227.065 117.350 ;
        RECT 272.090 117.180 272.260 117.350 ;
        RECT 272.450 117.180 272.620 117.350 ;
        RECT 272.810 117.180 272.980 117.350 ;
        RECT 273.170 117.180 273.340 117.350 ;
        RECT 273.530 117.180 273.700 117.350 ;
        RECT 273.890 117.180 274.060 117.350 ;
        RECT 147.205 116.130 147.375 116.300 ;
        RECT 147.565 116.130 147.735 116.300 ;
        RECT 147.925 116.130 148.095 116.300 ;
        RECT 148.285 116.130 148.455 116.300 ;
        RECT 148.645 116.130 148.815 116.300 ;
        RECT 149.005 116.130 149.175 116.300 ;
        RECT 194.200 116.130 194.370 116.300 ;
        RECT 194.560 116.130 194.730 116.300 ;
        RECT 194.920 116.130 195.090 116.300 ;
        RECT 195.280 116.130 195.450 116.300 ;
        RECT 195.640 116.130 195.810 116.300 ;
        RECT 196.000 116.130 196.170 116.300 ;
        RECT 199.265 116.100 201.235 116.630 ;
        RECT 220.260 116.100 222.230 116.630 ;
        RECT 225.095 116.350 225.265 116.520 ;
        RECT 225.455 116.350 225.625 116.520 ;
        RECT 225.815 116.350 225.985 116.520 ;
        RECT 226.175 116.350 226.345 116.520 ;
        RECT 226.535 116.350 226.705 116.520 ;
        RECT 226.895 116.350 227.065 116.520 ;
        RECT 272.090 116.350 272.260 116.520 ;
        RECT 272.450 116.350 272.620 116.520 ;
        RECT 272.810 116.350 272.980 116.520 ;
        RECT 273.170 116.350 273.340 116.520 ;
        RECT 273.530 116.350 273.700 116.520 ;
        RECT 273.890 116.350 274.060 116.520 ;
        RECT 147.205 115.300 147.375 115.470 ;
        RECT 147.565 115.300 147.735 115.470 ;
        RECT 147.925 115.300 148.095 115.470 ;
        RECT 148.285 115.300 148.455 115.470 ;
        RECT 148.645 115.300 148.815 115.470 ;
        RECT 149.005 115.300 149.175 115.470 ;
        RECT 194.200 115.300 194.370 115.470 ;
        RECT 194.560 115.300 194.730 115.470 ;
        RECT 194.920 115.300 195.090 115.470 ;
        RECT 195.280 115.300 195.450 115.470 ;
        RECT 195.640 115.300 195.810 115.470 ;
        RECT 196.000 115.300 196.170 115.470 ;
        RECT 199.265 114.930 201.235 115.460 ;
        RECT 220.260 114.930 222.230 115.460 ;
        RECT 225.095 115.520 225.265 115.690 ;
        RECT 225.455 115.520 225.625 115.690 ;
        RECT 225.815 115.520 225.985 115.690 ;
        RECT 226.175 115.520 226.345 115.690 ;
        RECT 226.535 115.520 226.705 115.690 ;
        RECT 226.895 115.520 227.065 115.690 ;
        RECT 272.090 115.520 272.260 115.690 ;
        RECT 272.450 115.520 272.620 115.690 ;
        RECT 272.810 115.520 272.980 115.690 ;
        RECT 273.170 115.520 273.340 115.690 ;
        RECT 273.530 115.520 273.700 115.690 ;
        RECT 273.890 115.520 274.060 115.690 ;
        RECT 147.205 114.470 147.375 114.640 ;
        RECT 147.565 114.470 147.735 114.640 ;
        RECT 147.925 114.470 148.095 114.640 ;
        RECT 148.285 114.470 148.455 114.640 ;
        RECT 148.645 114.470 148.815 114.640 ;
        RECT 149.005 114.470 149.175 114.640 ;
        RECT 194.200 114.470 194.370 114.640 ;
        RECT 194.560 114.470 194.730 114.640 ;
        RECT 194.920 114.470 195.090 114.640 ;
        RECT 195.280 114.470 195.450 114.640 ;
        RECT 195.640 114.470 195.810 114.640 ;
        RECT 196.000 114.470 196.170 114.640 ;
        RECT 225.095 114.690 225.265 114.860 ;
        RECT 225.455 114.690 225.625 114.860 ;
        RECT 225.815 114.690 225.985 114.860 ;
        RECT 226.175 114.690 226.345 114.860 ;
        RECT 226.535 114.690 226.705 114.860 ;
        RECT 226.895 114.690 227.065 114.860 ;
        RECT 272.090 114.690 272.260 114.860 ;
        RECT 272.450 114.690 272.620 114.860 ;
        RECT 272.810 114.690 272.980 114.860 ;
        RECT 273.170 114.690 273.340 114.860 ;
        RECT 273.530 114.690 273.700 114.860 ;
        RECT 273.890 114.690 274.060 114.860 ;
        RECT 147.205 113.640 147.375 113.810 ;
        RECT 147.565 113.640 147.735 113.810 ;
        RECT 147.925 113.640 148.095 113.810 ;
        RECT 148.285 113.640 148.455 113.810 ;
        RECT 148.645 113.640 148.815 113.810 ;
        RECT 149.005 113.640 149.175 113.810 ;
        RECT 194.200 113.640 194.370 113.810 ;
        RECT 194.560 113.640 194.730 113.810 ;
        RECT 194.920 113.640 195.090 113.810 ;
        RECT 195.280 113.640 195.450 113.810 ;
        RECT 195.640 113.640 195.810 113.810 ;
        RECT 196.000 113.640 196.170 113.810 ;
        RECT 199.265 113.760 201.235 114.290 ;
        RECT 220.260 113.760 222.230 114.290 ;
        RECT 225.095 113.860 225.265 114.030 ;
        RECT 225.455 113.860 225.625 114.030 ;
        RECT 225.815 113.860 225.985 114.030 ;
        RECT 226.175 113.860 226.345 114.030 ;
        RECT 226.535 113.860 226.705 114.030 ;
        RECT 226.895 113.860 227.065 114.030 ;
        RECT 272.090 113.860 272.260 114.030 ;
        RECT 272.450 113.860 272.620 114.030 ;
        RECT 272.810 113.860 272.980 114.030 ;
        RECT 273.170 113.860 273.340 114.030 ;
        RECT 273.530 113.860 273.700 114.030 ;
        RECT 273.890 113.860 274.060 114.030 ;
        RECT 147.205 112.810 147.375 112.980 ;
        RECT 147.565 112.810 147.735 112.980 ;
        RECT 147.925 112.810 148.095 112.980 ;
        RECT 148.285 112.810 148.455 112.980 ;
        RECT 148.645 112.810 148.815 112.980 ;
        RECT 149.005 112.810 149.175 112.980 ;
        RECT 194.200 112.810 194.370 112.980 ;
        RECT 194.560 112.810 194.730 112.980 ;
        RECT 194.920 112.810 195.090 112.980 ;
        RECT 195.280 112.810 195.450 112.980 ;
        RECT 195.640 112.810 195.810 112.980 ;
        RECT 196.000 112.810 196.170 112.980 ;
        RECT 199.265 112.590 201.235 113.120 ;
        RECT 220.260 112.590 222.230 113.120 ;
        RECT 225.095 113.030 225.265 113.200 ;
        RECT 225.455 113.030 225.625 113.200 ;
        RECT 225.815 113.030 225.985 113.200 ;
        RECT 226.175 113.030 226.345 113.200 ;
        RECT 226.535 113.030 226.705 113.200 ;
        RECT 226.895 113.030 227.065 113.200 ;
        RECT 272.090 113.030 272.260 113.200 ;
        RECT 272.450 113.030 272.620 113.200 ;
        RECT 272.810 113.030 272.980 113.200 ;
        RECT 273.170 113.030 273.340 113.200 ;
        RECT 273.530 113.030 273.700 113.200 ;
        RECT 273.890 113.030 274.060 113.200 ;
        RECT 147.205 111.980 147.375 112.150 ;
        RECT 147.565 111.980 147.735 112.150 ;
        RECT 147.925 111.980 148.095 112.150 ;
        RECT 148.285 111.980 148.455 112.150 ;
        RECT 148.645 111.980 148.815 112.150 ;
        RECT 149.005 111.980 149.175 112.150 ;
        RECT 194.200 111.980 194.370 112.150 ;
        RECT 194.560 111.980 194.730 112.150 ;
        RECT 194.920 111.980 195.090 112.150 ;
        RECT 195.280 111.980 195.450 112.150 ;
        RECT 195.640 111.980 195.810 112.150 ;
        RECT 196.000 111.980 196.170 112.150 ;
        RECT 225.095 112.200 225.265 112.370 ;
        RECT 225.455 112.200 225.625 112.370 ;
        RECT 225.815 112.200 225.985 112.370 ;
        RECT 226.175 112.200 226.345 112.370 ;
        RECT 226.535 112.200 226.705 112.370 ;
        RECT 226.895 112.200 227.065 112.370 ;
        RECT 272.090 112.200 272.260 112.370 ;
        RECT 272.450 112.200 272.620 112.370 ;
        RECT 272.810 112.200 272.980 112.370 ;
        RECT 273.170 112.200 273.340 112.370 ;
        RECT 273.530 112.200 273.700 112.370 ;
        RECT 273.890 112.200 274.060 112.370 ;
        RECT 199.265 111.420 201.235 111.950 ;
        RECT 147.205 111.150 147.375 111.320 ;
        RECT 147.565 111.150 147.735 111.320 ;
        RECT 147.925 111.150 148.095 111.320 ;
        RECT 148.285 111.150 148.455 111.320 ;
        RECT 148.645 111.150 148.815 111.320 ;
        RECT 149.005 111.150 149.175 111.320 ;
        RECT 220.260 111.420 222.230 111.950 ;
        RECT 225.095 111.370 225.265 111.540 ;
        RECT 225.455 111.370 225.625 111.540 ;
        RECT 225.815 111.370 225.985 111.540 ;
        RECT 226.175 111.370 226.345 111.540 ;
        RECT 226.535 111.370 226.705 111.540 ;
        RECT 226.895 111.370 227.065 111.540 ;
        RECT 194.200 111.150 194.370 111.320 ;
        RECT 194.560 111.150 194.730 111.320 ;
        RECT 194.920 111.150 195.090 111.320 ;
        RECT 195.280 111.150 195.450 111.320 ;
        RECT 195.640 111.150 195.810 111.320 ;
        RECT 196.000 111.150 196.170 111.320 ;
        RECT 272.090 111.370 272.260 111.540 ;
        RECT 272.450 111.370 272.620 111.540 ;
        RECT 272.810 111.370 272.980 111.540 ;
        RECT 273.170 111.370 273.340 111.540 ;
        RECT 273.530 111.370 273.700 111.540 ;
        RECT 273.890 111.370 274.060 111.540 ;
        RECT 147.205 110.320 147.375 110.490 ;
        RECT 147.565 110.320 147.735 110.490 ;
        RECT 147.925 110.320 148.095 110.490 ;
        RECT 148.285 110.320 148.455 110.490 ;
        RECT 148.645 110.320 148.815 110.490 ;
        RECT 149.005 110.320 149.175 110.490 ;
        RECT 194.200 110.320 194.370 110.490 ;
        RECT 194.560 110.320 194.730 110.490 ;
        RECT 194.920 110.320 195.090 110.490 ;
        RECT 195.280 110.320 195.450 110.490 ;
        RECT 195.640 110.320 195.810 110.490 ;
        RECT 196.000 110.320 196.170 110.490 ;
        RECT 199.265 110.250 201.235 110.780 ;
        RECT 220.260 110.250 222.230 110.780 ;
        RECT 225.095 110.540 225.265 110.710 ;
        RECT 225.455 110.540 225.625 110.710 ;
        RECT 225.815 110.540 225.985 110.710 ;
        RECT 226.175 110.540 226.345 110.710 ;
        RECT 226.535 110.540 226.705 110.710 ;
        RECT 226.895 110.540 227.065 110.710 ;
        RECT 272.090 110.540 272.260 110.710 ;
        RECT 272.450 110.540 272.620 110.710 ;
        RECT 272.810 110.540 272.980 110.710 ;
        RECT 273.170 110.540 273.340 110.710 ;
        RECT 273.530 110.540 273.700 110.710 ;
        RECT 273.890 110.540 274.060 110.710 ;
        RECT 147.205 109.490 147.375 109.660 ;
        RECT 147.565 109.490 147.735 109.660 ;
        RECT 147.925 109.490 148.095 109.660 ;
        RECT 148.285 109.490 148.455 109.660 ;
        RECT 148.645 109.490 148.815 109.660 ;
        RECT 149.005 109.490 149.175 109.660 ;
        RECT 225.095 109.710 225.265 109.880 ;
        RECT 225.455 109.710 225.625 109.880 ;
        RECT 225.815 109.710 225.985 109.880 ;
        RECT 226.175 109.710 226.345 109.880 ;
        RECT 226.535 109.710 226.705 109.880 ;
        RECT 226.895 109.710 227.065 109.880 ;
        RECT 194.200 109.490 194.370 109.660 ;
        RECT 194.560 109.490 194.730 109.660 ;
        RECT 194.920 109.490 195.090 109.660 ;
        RECT 195.280 109.490 195.450 109.660 ;
        RECT 195.640 109.490 195.810 109.660 ;
        RECT 196.000 109.490 196.170 109.660 ;
        RECT 199.265 109.080 201.235 109.610 ;
        RECT 272.090 109.710 272.260 109.880 ;
        RECT 272.450 109.710 272.620 109.880 ;
        RECT 272.810 109.710 272.980 109.880 ;
        RECT 273.170 109.710 273.340 109.880 ;
        RECT 273.530 109.710 273.700 109.880 ;
        RECT 273.890 109.710 274.060 109.880 ;
        RECT 220.260 109.080 222.230 109.610 ;
        RECT 147.205 108.660 147.375 108.830 ;
        RECT 147.565 108.660 147.735 108.830 ;
        RECT 147.925 108.660 148.095 108.830 ;
        RECT 148.285 108.660 148.455 108.830 ;
        RECT 148.645 108.660 148.815 108.830 ;
        RECT 149.005 108.660 149.175 108.830 ;
        RECT 194.200 108.660 194.370 108.830 ;
        RECT 194.560 108.660 194.730 108.830 ;
        RECT 194.920 108.660 195.090 108.830 ;
        RECT 195.280 108.660 195.450 108.830 ;
        RECT 195.640 108.660 195.810 108.830 ;
        RECT 196.000 108.660 196.170 108.830 ;
        RECT 225.095 108.880 225.265 109.050 ;
        RECT 225.455 108.880 225.625 109.050 ;
        RECT 225.815 108.880 225.985 109.050 ;
        RECT 226.175 108.880 226.345 109.050 ;
        RECT 226.535 108.880 226.705 109.050 ;
        RECT 226.895 108.880 227.065 109.050 ;
        RECT 272.090 108.880 272.260 109.050 ;
        RECT 272.450 108.880 272.620 109.050 ;
        RECT 272.810 108.880 272.980 109.050 ;
        RECT 273.170 108.880 273.340 109.050 ;
        RECT 273.530 108.880 273.700 109.050 ;
        RECT 273.890 108.880 274.060 109.050 ;
        RECT 147.205 107.830 147.375 108.000 ;
        RECT 147.565 107.830 147.735 108.000 ;
        RECT 147.925 107.830 148.095 108.000 ;
        RECT 148.285 107.830 148.455 108.000 ;
        RECT 148.645 107.830 148.815 108.000 ;
        RECT 149.005 107.830 149.175 108.000 ;
        RECT 194.200 107.830 194.370 108.000 ;
        RECT 194.560 107.830 194.730 108.000 ;
        RECT 194.920 107.830 195.090 108.000 ;
        RECT 195.280 107.830 195.450 108.000 ;
        RECT 195.640 107.830 195.810 108.000 ;
        RECT 196.000 107.830 196.170 108.000 ;
        RECT 199.265 107.910 201.235 108.440 ;
        RECT 220.260 107.910 222.230 108.440 ;
        RECT 225.095 108.050 225.265 108.220 ;
        RECT 225.455 108.050 225.625 108.220 ;
        RECT 225.815 108.050 225.985 108.220 ;
        RECT 226.175 108.050 226.345 108.220 ;
        RECT 226.535 108.050 226.705 108.220 ;
        RECT 226.895 108.050 227.065 108.220 ;
        RECT 272.090 108.050 272.260 108.220 ;
        RECT 272.450 108.050 272.620 108.220 ;
        RECT 272.810 108.050 272.980 108.220 ;
        RECT 273.170 108.050 273.340 108.220 ;
        RECT 273.530 108.050 273.700 108.220 ;
        RECT 273.890 108.050 274.060 108.220 ;
        RECT 147.205 107.000 147.375 107.170 ;
        RECT 147.565 107.000 147.735 107.170 ;
        RECT 147.925 107.000 148.095 107.170 ;
        RECT 148.285 107.000 148.455 107.170 ;
        RECT 148.645 107.000 148.815 107.170 ;
        RECT 149.005 107.000 149.175 107.170 ;
        RECT 194.200 107.000 194.370 107.170 ;
        RECT 194.560 107.000 194.730 107.170 ;
        RECT 194.920 107.000 195.090 107.170 ;
        RECT 195.280 107.000 195.450 107.170 ;
        RECT 195.640 107.000 195.810 107.170 ;
        RECT 196.000 107.000 196.170 107.170 ;
        RECT 199.265 106.740 201.235 107.270 ;
        RECT 220.260 106.740 222.230 107.270 ;
        RECT 225.095 107.220 225.265 107.390 ;
        RECT 225.455 107.220 225.625 107.390 ;
        RECT 225.815 107.220 225.985 107.390 ;
        RECT 226.175 107.220 226.345 107.390 ;
        RECT 226.535 107.220 226.705 107.390 ;
        RECT 226.895 107.220 227.065 107.390 ;
        RECT 272.090 107.220 272.260 107.390 ;
        RECT 272.450 107.220 272.620 107.390 ;
        RECT 272.810 107.220 272.980 107.390 ;
        RECT 273.170 107.220 273.340 107.390 ;
        RECT 273.530 107.220 273.700 107.390 ;
        RECT 273.890 107.220 274.060 107.390 ;
        RECT 147.205 106.170 147.375 106.340 ;
        RECT 147.565 106.170 147.735 106.340 ;
        RECT 147.925 106.170 148.095 106.340 ;
        RECT 148.285 106.170 148.455 106.340 ;
        RECT 148.645 106.170 148.815 106.340 ;
        RECT 149.005 106.170 149.175 106.340 ;
        RECT 194.200 106.170 194.370 106.340 ;
        RECT 194.560 106.170 194.730 106.340 ;
        RECT 194.920 106.170 195.090 106.340 ;
        RECT 195.280 106.170 195.450 106.340 ;
        RECT 195.640 106.170 195.810 106.340 ;
        RECT 196.000 106.170 196.170 106.340 ;
        RECT 225.095 106.390 225.265 106.560 ;
        RECT 225.455 106.390 225.625 106.560 ;
        RECT 225.815 106.390 225.985 106.560 ;
        RECT 226.175 106.390 226.345 106.560 ;
        RECT 226.535 106.390 226.705 106.560 ;
        RECT 226.895 106.390 227.065 106.560 ;
        RECT 272.090 106.390 272.260 106.560 ;
        RECT 272.450 106.390 272.620 106.560 ;
        RECT 272.810 106.390 272.980 106.560 ;
        RECT 273.170 106.390 273.340 106.560 ;
        RECT 273.530 106.390 273.700 106.560 ;
        RECT 273.890 106.390 274.060 106.560 ;
        RECT 147.205 105.340 147.375 105.510 ;
        RECT 147.565 105.340 147.735 105.510 ;
        RECT 147.925 105.340 148.095 105.510 ;
        RECT 148.285 105.340 148.455 105.510 ;
        RECT 148.645 105.340 148.815 105.510 ;
        RECT 149.005 105.340 149.175 105.510 ;
        RECT 194.200 105.340 194.370 105.510 ;
        RECT 194.560 105.340 194.730 105.510 ;
        RECT 194.920 105.340 195.090 105.510 ;
        RECT 195.280 105.340 195.450 105.510 ;
        RECT 195.640 105.340 195.810 105.510 ;
        RECT 196.000 105.340 196.170 105.510 ;
        RECT 199.265 105.570 201.235 106.100 ;
        RECT 220.260 105.570 222.230 106.100 ;
        RECT 225.095 105.560 225.265 105.730 ;
        RECT 225.455 105.560 225.625 105.730 ;
        RECT 225.815 105.560 225.985 105.730 ;
        RECT 226.175 105.560 226.345 105.730 ;
        RECT 226.535 105.560 226.705 105.730 ;
        RECT 226.895 105.560 227.065 105.730 ;
        RECT 272.090 105.560 272.260 105.730 ;
        RECT 272.450 105.560 272.620 105.730 ;
        RECT 272.810 105.560 272.980 105.730 ;
        RECT 273.170 105.560 273.340 105.730 ;
        RECT 273.530 105.560 273.700 105.730 ;
        RECT 273.890 105.560 274.060 105.730 ;
        RECT 147.205 104.510 147.375 104.680 ;
        RECT 147.565 104.510 147.735 104.680 ;
        RECT 147.925 104.510 148.095 104.680 ;
        RECT 148.285 104.510 148.455 104.680 ;
        RECT 148.645 104.510 148.815 104.680 ;
        RECT 149.005 104.510 149.175 104.680 ;
        RECT 194.200 104.510 194.370 104.680 ;
        RECT 194.560 104.510 194.730 104.680 ;
        RECT 194.920 104.510 195.090 104.680 ;
        RECT 195.280 104.510 195.450 104.680 ;
        RECT 195.640 104.510 195.810 104.680 ;
        RECT 196.000 104.510 196.170 104.680 ;
        RECT 199.265 104.400 201.235 104.930 ;
        RECT 220.260 104.400 222.230 104.930 ;
        RECT 225.095 104.730 225.265 104.900 ;
        RECT 225.455 104.730 225.625 104.900 ;
        RECT 225.815 104.730 225.985 104.900 ;
        RECT 226.175 104.730 226.345 104.900 ;
        RECT 226.535 104.730 226.705 104.900 ;
        RECT 226.895 104.730 227.065 104.900 ;
        RECT 272.090 104.730 272.260 104.900 ;
        RECT 272.450 104.730 272.620 104.900 ;
        RECT 272.810 104.730 272.980 104.900 ;
        RECT 273.170 104.730 273.340 104.900 ;
        RECT 273.530 104.730 273.700 104.900 ;
        RECT 273.890 104.730 274.060 104.900 ;
        RECT 147.205 103.680 147.375 103.850 ;
        RECT 147.565 103.680 147.735 103.850 ;
        RECT 147.925 103.680 148.095 103.850 ;
        RECT 148.285 103.680 148.455 103.850 ;
        RECT 148.645 103.680 148.815 103.850 ;
        RECT 149.005 103.680 149.175 103.850 ;
        RECT 194.200 103.680 194.370 103.850 ;
        RECT 194.560 103.680 194.730 103.850 ;
        RECT 194.920 103.680 195.090 103.850 ;
        RECT 195.280 103.680 195.450 103.850 ;
        RECT 195.640 103.680 195.810 103.850 ;
        RECT 196.000 103.680 196.170 103.850 ;
        RECT 225.095 103.900 225.265 104.070 ;
        RECT 225.455 103.900 225.625 104.070 ;
        RECT 225.815 103.900 225.985 104.070 ;
        RECT 226.175 103.900 226.345 104.070 ;
        RECT 226.535 103.900 226.705 104.070 ;
        RECT 226.895 103.900 227.065 104.070 ;
        RECT 199.265 103.230 201.235 103.760 ;
        RECT 272.090 103.900 272.260 104.070 ;
        RECT 272.450 103.900 272.620 104.070 ;
        RECT 272.810 103.900 272.980 104.070 ;
        RECT 273.170 103.900 273.340 104.070 ;
        RECT 273.530 103.900 273.700 104.070 ;
        RECT 273.890 103.900 274.060 104.070 ;
        RECT 220.260 103.230 222.230 103.760 ;
        RECT 147.205 102.850 147.375 103.020 ;
        RECT 147.565 102.850 147.735 103.020 ;
        RECT 147.925 102.850 148.095 103.020 ;
        RECT 148.285 102.850 148.455 103.020 ;
        RECT 148.645 102.850 148.815 103.020 ;
        RECT 149.005 102.850 149.175 103.020 ;
        RECT 194.200 102.850 194.370 103.020 ;
        RECT 194.560 102.850 194.730 103.020 ;
        RECT 194.920 102.850 195.090 103.020 ;
        RECT 195.280 102.850 195.450 103.020 ;
        RECT 195.640 102.850 195.810 103.020 ;
        RECT 196.000 102.850 196.170 103.020 ;
        RECT 225.095 103.070 225.265 103.240 ;
        RECT 225.455 103.070 225.625 103.240 ;
        RECT 225.815 103.070 225.985 103.240 ;
        RECT 226.175 103.070 226.345 103.240 ;
        RECT 226.535 103.070 226.705 103.240 ;
        RECT 226.895 103.070 227.065 103.240 ;
        RECT 272.090 103.070 272.260 103.240 ;
        RECT 272.450 103.070 272.620 103.240 ;
        RECT 272.810 103.070 272.980 103.240 ;
        RECT 273.170 103.070 273.340 103.240 ;
        RECT 273.530 103.070 273.700 103.240 ;
        RECT 273.890 103.070 274.060 103.240 ;
        RECT 147.205 102.020 147.375 102.190 ;
        RECT 147.565 102.020 147.735 102.190 ;
        RECT 147.925 102.020 148.095 102.190 ;
        RECT 148.285 102.020 148.455 102.190 ;
        RECT 148.645 102.020 148.815 102.190 ;
        RECT 149.005 102.020 149.175 102.190 ;
        RECT 194.200 102.020 194.370 102.190 ;
        RECT 194.560 102.020 194.730 102.190 ;
        RECT 194.920 102.020 195.090 102.190 ;
        RECT 195.280 102.020 195.450 102.190 ;
        RECT 195.640 102.020 195.810 102.190 ;
        RECT 196.000 102.020 196.170 102.190 ;
        RECT 225.095 102.240 225.265 102.410 ;
        RECT 225.455 102.240 225.625 102.410 ;
        RECT 225.815 102.240 225.985 102.410 ;
        RECT 226.175 102.240 226.345 102.410 ;
        RECT 226.535 102.240 226.705 102.410 ;
        RECT 226.895 102.240 227.065 102.410 ;
        RECT 272.090 102.240 272.260 102.410 ;
        RECT 272.450 102.240 272.620 102.410 ;
        RECT 272.810 102.240 272.980 102.410 ;
        RECT 273.170 102.240 273.340 102.410 ;
        RECT 273.530 102.240 273.700 102.410 ;
        RECT 273.890 102.240 274.060 102.410 ;
        RECT 147.205 101.190 147.375 101.360 ;
        RECT 147.565 101.190 147.735 101.360 ;
        RECT 147.925 101.190 148.095 101.360 ;
        RECT 148.285 101.190 148.455 101.360 ;
        RECT 148.645 101.190 148.815 101.360 ;
        RECT 149.005 101.190 149.175 101.360 ;
        RECT 194.200 101.190 194.370 101.360 ;
        RECT 194.560 101.190 194.730 101.360 ;
        RECT 194.920 101.190 195.090 101.360 ;
        RECT 195.280 101.190 195.450 101.360 ;
        RECT 195.640 101.190 195.810 101.360 ;
        RECT 196.000 101.190 196.170 101.360 ;
        RECT 225.095 101.410 225.265 101.580 ;
        RECT 225.455 101.410 225.625 101.580 ;
        RECT 225.815 101.410 225.985 101.580 ;
        RECT 226.175 101.410 226.345 101.580 ;
        RECT 226.535 101.410 226.705 101.580 ;
        RECT 226.895 101.410 227.065 101.580 ;
        RECT 272.090 101.410 272.260 101.580 ;
        RECT 272.450 101.410 272.620 101.580 ;
        RECT 272.810 101.410 272.980 101.580 ;
        RECT 273.170 101.410 273.340 101.580 ;
        RECT 273.530 101.410 273.700 101.580 ;
        RECT 273.890 101.410 274.060 101.580 ;
        RECT 147.205 100.360 147.375 100.530 ;
        RECT 147.565 100.360 147.735 100.530 ;
        RECT 147.925 100.360 148.095 100.530 ;
        RECT 148.285 100.360 148.455 100.530 ;
        RECT 148.645 100.360 148.815 100.530 ;
        RECT 149.005 100.360 149.175 100.530 ;
        RECT 194.200 100.360 194.370 100.530 ;
        RECT 194.560 100.360 194.730 100.530 ;
        RECT 194.920 100.360 195.090 100.530 ;
        RECT 195.280 100.360 195.450 100.530 ;
        RECT 195.640 100.360 195.810 100.530 ;
        RECT 196.000 100.360 196.170 100.530 ;
        RECT 225.095 100.580 225.265 100.750 ;
        RECT 225.455 100.580 225.625 100.750 ;
        RECT 225.815 100.580 225.985 100.750 ;
        RECT 226.175 100.580 226.345 100.750 ;
        RECT 226.535 100.580 226.705 100.750 ;
        RECT 226.895 100.580 227.065 100.750 ;
        RECT 272.090 100.580 272.260 100.750 ;
        RECT 272.450 100.580 272.620 100.750 ;
        RECT 272.810 100.580 272.980 100.750 ;
        RECT 273.170 100.580 273.340 100.750 ;
        RECT 273.530 100.580 273.700 100.750 ;
        RECT 273.890 100.580 274.060 100.750 ;
        RECT 147.205 99.530 147.375 99.700 ;
        RECT 147.565 99.530 147.735 99.700 ;
        RECT 147.925 99.530 148.095 99.700 ;
        RECT 148.285 99.530 148.455 99.700 ;
        RECT 148.645 99.530 148.815 99.700 ;
        RECT 149.005 99.530 149.175 99.700 ;
        RECT 194.200 99.530 194.370 99.700 ;
        RECT 194.560 99.530 194.730 99.700 ;
        RECT 194.920 99.530 195.090 99.700 ;
        RECT 195.280 99.530 195.450 99.700 ;
        RECT 195.640 99.530 195.810 99.700 ;
        RECT 196.000 99.530 196.170 99.700 ;
        RECT 225.095 99.750 225.265 99.920 ;
        RECT 225.455 99.750 225.625 99.920 ;
        RECT 225.815 99.750 225.985 99.920 ;
        RECT 226.175 99.750 226.345 99.920 ;
        RECT 226.535 99.750 226.705 99.920 ;
        RECT 226.895 99.750 227.065 99.920 ;
        RECT 272.090 99.750 272.260 99.920 ;
        RECT 272.450 99.750 272.620 99.920 ;
        RECT 272.810 99.750 272.980 99.920 ;
        RECT 273.170 99.750 273.340 99.920 ;
        RECT 273.530 99.750 273.700 99.920 ;
        RECT 273.890 99.750 274.060 99.920 ;
        RECT 212.370 99.180 212.540 99.350 ;
        RECT 215.060 99.180 215.230 99.350 ;
        RECT 147.205 98.700 147.375 98.870 ;
        RECT 147.565 98.700 147.735 98.870 ;
        RECT 147.925 98.700 148.095 98.870 ;
        RECT 148.285 98.700 148.455 98.870 ;
        RECT 148.645 98.700 148.815 98.870 ;
        RECT 149.005 98.700 149.175 98.870 ;
        RECT 194.200 98.700 194.370 98.870 ;
        RECT 194.560 98.700 194.730 98.870 ;
        RECT 194.920 98.700 195.090 98.870 ;
        RECT 195.280 98.700 195.450 98.870 ;
        RECT 195.640 98.700 195.810 98.870 ;
        RECT 196.000 98.700 196.170 98.870 ;
        RECT 208.080 98.700 208.250 98.870 ;
        RECT 211.885 98.785 212.055 98.955 ;
        RECT 215.545 98.785 215.715 98.955 ;
        RECT 225.095 98.920 225.265 99.090 ;
        RECT 225.455 98.920 225.625 99.090 ;
        RECT 225.815 98.920 225.985 99.090 ;
        RECT 226.175 98.920 226.345 99.090 ;
        RECT 226.535 98.920 226.705 99.090 ;
        RECT 226.895 98.920 227.065 99.090 ;
        RECT 272.090 98.920 272.260 99.090 ;
        RECT 272.450 98.920 272.620 99.090 ;
        RECT 272.810 98.920 272.980 99.090 ;
        RECT 273.170 98.920 273.340 99.090 ;
        RECT 273.530 98.920 273.700 99.090 ;
        RECT 273.890 98.920 274.060 99.090 ;
        RECT 208.610 98.305 208.780 98.475 ;
        RECT 212.370 98.390 212.540 98.560 ;
        RECT 147.205 97.870 147.375 98.040 ;
        RECT 147.565 97.870 147.735 98.040 ;
        RECT 147.925 97.870 148.095 98.040 ;
        RECT 148.285 97.870 148.455 98.040 ;
        RECT 148.645 97.870 148.815 98.040 ;
        RECT 149.005 97.870 149.175 98.040 ;
        RECT 194.200 97.870 194.370 98.040 ;
        RECT 194.560 97.870 194.730 98.040 ;
        RECT 194.920 97.870 195.090 98.040 ;
        RECT 195.280 97.870 195.450 98.040 ;
        RECT 195.640 97.870 195.810 98.040 ;
        RECT 196.000 97.870 196.170 98.040 ;
        RECT 225.095 98.090 225.265 98.260 ;
        RECT 225.455 98.090 225.625 98.260 ;
        RECT 225.815 98.090 225.985 98.260 ;
        RECT 226.175 98.090 226.345 98.260 ;
        RECT 226.535 98.090 226.705 98.260 ;
        RECT 226.895 98.090 227.065 98.260 ;
        RECT 272.090 98.090 272.260 98.260 ;
        RECT 272.450 98.090 272.620 98.260 ;
        RECT 272.810 98.090 272.980 98.260 ;
        RECT 273.170 98.090 273.340 98.260 ;
        RECT 273.530 98.090 273.700 98.260 ;
        RECT 273.890 98.090 274.060 98.260 ;
        RECT 147.205 97.040 147.375 97.210 ;
        RECT 147.565 97.040 147.735 97.210 ;
        RECT 147.925 97.040 148.095 97.210 ;
        RECT 148.285 97.040 148.455 97.210 ;
        RECT 148.645 97.040 148.815 97.210 ;
        RECT 149.005 97.040 149.175 97.210 ;
        RECT 194.200 97.040 194.370 97.210 ;
        RECT 194.560 97.040 194.730 97.210 ;
        RECT 194.920 97.040 195.090 97.210 ;
        RECT 195.280 97.040 195.450 97.210 ;
        RECT 195.640 97.040 195.810 97.210 ;
        RECT 196.000 97.040 196.170 97.210 ;
        RECT 225.095 97.260 225.265 97.430 ;
        RECT 225.455 97.260 225.625 97.430 ;
        RECT 225.815 97.260 225.985 97.430 ;
        RECT 226.175 97.260 226.345 97.430 ;
        RECT 226.535 97.260 226.705 97.430 ;
        RECT 226.895 97.260 227.065 97.430 ;
        RECT 272.090 97.260 272.260 97.430 ;
        RECT 272.450 97.260 272.620 97.430 ;
        RECT 272.810 97.260 272.980 97.430 ;
        RECT 273.170 97.260 273.340 97.430 ;
        RECT 273.530 97.260 273.700 97.430 ;
        RECT 273.890 97.260 274.060 97.430 ;
        RECT 147.205 96.210 147.375 96.380 ;
        RECT 147.565 96.210 147.735 96.380 ;
        RECT 147.925 96.210 148.095 96.380 ;
        RECT 148.285 96.210 148.455 96.380 ;
        RECT 148.645 96.210 148.815 96.380 ;
        RECT 149.005 96.210 149.175 96.380 ;
        RECT 212.370 96.400 212.540 96.570 ;
        RECT 215.060 96.400 215.230 96.570 ;
        RECT 225.095 96.430 225.265 96.600 ;
        RECT 225.455 96.430 225.625 96.600 ;
        RECT 225.815 96.430 225.985 96.600 ;
        RECT 226.175 96.430 226.345 96.600 ;
        RECT 226.535 96.430 226.705 96.600 ;
        RECT 226.895 96.430 227.065 96.600 ;
        RECT 194.200 96.210 194.370 96.380 ;
        RECT 194.560 96.210 194.730 96.380 ;
        RECT 194.920 96.210 195.090 96.380 ;
        RECT 195.280 96.210 195.450 96.380 ;
        RECT 195.640 96.210 195.810 96.380 ;
        RECT 196.000 96.210 196.170 96.380 ;
        RECT 272.090 96.430 272.260 96.600 ;
        RECT 272.450 96.430 272.620 96.600 ;
        RECT 272.810 96.430 272.980 96.600 ;
        RECT 273.170 96.430 273.340 96.600 ;
        RECT 273.530 96.430 273.700 96.600 ;
        RECT 273.890 96.430 274.060 96.600 ;
        RECT 211.885 96.005 212.055 96.175 ;
        RECT 215.545 96.005 215.715 96.175 ;
        RECT 147.205 95.380 147.375 95.550 ;
        RECT 147.565 95.380 147.735 95.550 ;
        RECT 147.925 95.380 148.095 95.550 ;
        RECT 148.285 95.380 148.455 95.550 ;
        RECT 148.645 95.380 148.815 95.550 ;
        RECT 149.005 95.380 149.175 95.550 ;
        RECT 208.080 95.620 208.250 95.790 ;
        RECT 212.370 95.610 212.540 95.780 ;
        RECT 225.095 95.600 225.265 95.770 ;
        RECT 225.455 95.600 225.625 95.770 ;
        RECT 225.815 95.600 225.985 95.770 ;
        RECT 226.175 95.600 226.345 95.770 ;
        RECT 226.535 95.600 226.705 95.770 ;
        RECT 226.895 95.600 227.065 95.770 ;
        RECT 194.200 95.380 194.370 95.550 ;
        RECT 194.560 95.380 194.730 95.550 ;
        RECT 194.920 95.380 195.090 95.550 ;
        RECT 195.280 95.380 195.450 95.550 ;
        RECT 195.640 95.380 195.810 95.550 ;
        RECT 196.000 95.380 196.170 95.550 ;
        RECT 204.520 95.225 204.690 95.395 ;
        RECT 272.090 95.600 272.260 95.770 ;
        RECT 272.450 95.600 272.620 95.770 ;
        RECT 272.810 95.600 272.980 95.770 ;
        RECT 273.170 95.600 273.340 95.770 ;
        RECT 273.530 95.600 273.700 95.770 ;
        RECT 273.890 95.600 274.060 95.770 ;
        RECT 208.610 95.225 208.780 95.395 ;
        RECT 205.050 94.830 205.220 95.000 ;
        RECT 208.080 94.830 208.250 95.000 ;
        RECT 147.205 94.550 147.375 94.720 ;
        RECT 147.565 94.550 147.735 94.720 ;
        RECT 147.925 94.550 148.095 94.720 ;
        RECT 148.285 94.550 148.455 94.720 ;
        RECT 148.645 94.550 148.815 94.720 ;
        RECT 149.005 94.550 149.175 94.720 ;
        RECT 194.200 94.550 194.370 94.720 ;
        RECT 194.560 94.550 194.730 94.720 ;
        RECT 194.920 94.550 195.090 94.720 ;
        RECT 195.280 94.550 195.450 94.720 ;
        RECT 195.640 94.550 195.810 94.720 ;
        RECT 196.000 94.550 196.170 94.720 ;
        RECT 225.095 94.770 225.265 94.940 ;
        RECT 225.455 94.770 225.625 94.940 ;
        RECT 225.815 94.770 225.985 94.940 ;
        RECT 226.175 94.770 226.345 94.940 ;
        RECT 226.535 94.770 226.705 94.940 ;
        RECT 226.895 94.770 227.065 94.940 ;
        RECT 272.090 94.770 272.260 94.940 ;
        RECT 272.450 94.770 272.620 94.940 ;
        RECT 272.810 94.770 272.980 94.940 ;
        RECT 273.170 94.770 273.340 94.940 ;
        RECT 273.530 94.770 273.700 94.940 ;
        RECT 273.890 94.770 274.060 94.940 ;
        RECT 147.205 93.720 147.375 93.890 ;
        RECT 147.565 93.720 147.735 93.890 ;
        RECT 147.925 93.720 148.095 93.890 ;
        RECT 148.285 93.720 148.455 93.890 ;
        RECT 148.645 93.720 148.815 93.890 ;
        RECT 149.005 93.720 149.175 93.890 ;
        RECT 194.200 93.720 194.370 93.890 ;
        RECT 194.560 93.720 194.730 93.890 ;
        RECT 194.920 93.720 195.090 93.890 ;
        RECT 195.280 93.720 195.450 93.890 ;
        RECT 195.640 93.720 195.810 93.890 ;
        RECT 196.000 93.720 196.170 93.890 ;
        RECT 225.095 93.940 225.265 94.110 ;
        RECT 225.455 93.940 225.625 94.110 ;
        RECT 225.815 93.940 225.985 94.110 ;
        RECT 226.175 93.940 226.345 94.110 ;
        RECT 226.535 93.940 226.705 94.110 ;
        RECT 226.895 93.940 227.065 94.110 ;
        RECT 272.090 93.940 272.260 94.110 ;
        RECT 272.450 93.940 272.620 94.110 ;
        RECT 272.810 93.940 272.980 94.110 ;
        RECT 273.170 93.940 273.340 94.110 ;
        RECT 273.530 93.940 273.700 94.110 ;
        RECT 273.890 93.940 274.060 94.110 ;
        RECT 212.370 93.620 212.540 93.790 ;
        RECT 215.060 93.620 215.230 93.790 ;
        RECT 218.690 93.610 218.860 93.780 ;
        RECT 211.885 93.225 212.055 93.395 ;
        RECT 147.205 92.890 147.375 93.060 ;
        RECT 147.565 92.890 147.735 93.060 ;
        RECT 147.925 92.890 148.095 93.060 ;
        RECT 148.285 92.890 148.455 93.060 ;
        RECT 148.645 92.890 148.815 93.060 ;
        RECT 149.005 92.890 149.175 93.060 ;
        RECT 215.545 93.225 215.715 93.395 ;
        RECT 219.175 93.215 219.345 93.385 ;
        RECT 194.200 92.890 194.370 93.060 ;
        RECT 194.560 92.890 194.730 93.060 ;
        RECT 194.920 92.890 195.090 93.060 ;
        RECT 195.280 92.890 195.450 93.060 ;
        RECT 195.640 92.890 195.810 93.060 ;
        RECT 196.000 92.890 196.170 93.060 ;
        RECT 225.095 93.110 225.265 93.280 ;
        RECT 225.455 93.110 225.625 93.280 ;
        RECT 225.815 93.110 225.985 93.280 ;
        RECT 226.175 93.110 226.345 93.280 ;
        RECT 226.535 93.110 226.705 93.280 ;
        RECT 226.895 93.110 227.065 93.280 ;
        RECT 272.090 93.110 272.260 93.280 ;
        RECT 272.450 93.110 272.620 93.280 ;
        RECT 272.810 93.110 272.980 93.280 ;
        RECT 273.170 93.110 273.340 93.280 ;
        RECT 273.530 93.110 273.700 93.280 ;
        RECT 273.890 93.110 274.060 93.280 ;
        RECT 212.370 92.830 212.540 93.000 ;
        RECT 208.080 92.540 208.250 92.710 ;
        RECT 147.205 92.060 147.375 92.230 ;
        RECT 147.565 92.060 147.735 92.230 ;
        RECT 147.925 92.060 148.095 92.230 ;
        RECT 148.285 92.060 148.455 92.230 ;
        RECT 148.645 92.060 148.815 92.230 ;
        RECT 149.005 92.060 149.175 92.230 ;
        RECT 194.200 92.060 194.370 92.230 ;
        RECT 194.560 92.060 194.730 92.230 ;
        RECT 194.920 92.060 195.090 92.230 ;
        RECT 195.280 92.060 195.450 92.230 ;
        RECT 195.640 92.060 195.810 92.230 ;
        RECT 196.000 92.060 196.170 92.230 ;
        RECT 204.520 92.145 204.690 92.315 ;
        RECT 208.610 92.145 208.780 92.315 ;
        RECT 225.095 92.280 225.265 92.450 ;
        RECT 225.455 92.280 225.625 92.450 ;
        RECT 225.815 92.280 225.985 92.450 ;
        RECT 226.175 92.280 226.345 92.450 ;
        RECT 226.535 92.280 226.705 92.450 ;
        RECT 226.895 92.280 227.065 92.450 ;
        RECT 272.090 92.280 272.260 92.450 ;
        RECT 272.450 92.280 272.620 92.450 ;
        RECT 272.810 92.280 272.980 92.450 ;
        RECT 273.170 92.280 273.340 92.450 ;
        RECT 273.530 92.280 273.700 92.450 ;
        RECT 273.890 92.280 274.060 92.450 ;
        RECT 205.050 91.750 205.220 91.920 ;
        RECT 208.080 91.750 208.250 91.920 ;
        RECT 147.205 91.230 147.375 91.400 ;
        RECT 147.565 91.230 147.735 91.400 ;
        RECT 147.925 91.230 148.095 91.400 ;
        RECT 148.285 91.230 148.455 91.400 ;
        RECT 148.645 91.230 148.815 91.400 ;
        RECT 149.005 91.230 149.175 91.400 ;
        RECT 194.200 91.230 194.370 91.400 ;
        RECT 194.560 91.230 194.730 91.400 ;
        RECT 194.920 91.230 195.090 91.400 ;
        RECT 195.280 91.230 195.450 91.400 ;
        RECT 195.640 91.230 195.810 91.400 ;
        RECT 196.000 91.230 196.170 91.400 ;
        RECT 225.095 91.450 225.265 91.620 ;
        RECT 225.455 91.450 225.625 91.620 ;
        RECT 225.815 91.450 225.985 91.620 ;
        RECT 226.175 91.450 226.345 91.620 ;
        RECT 226.535 91.450 226.705 91.620 ;
        RECT 226.895 91.450 227.065 91.620 ;
        RECT 272.090 91.450 272.260 91.620 ;
        RECT 272.450 91.450 272.620 91.620 ;
        RECT 272.810 91.450 272.980 91.620 ;
        RECT 273.170 91.450 273.340 91.620 ;
        RECT 273.530 91.450 273.700 91.620 ;
        RECT 273.890 91.450 274.060 91.620 ;
        RECT 212.370 90.840 212.540 91.010 ;
        RECT 215.060 90.840 215.230 91.010 ;
        RECT 147.205 90.400 147.375 90.570 ;
        RECT 147.565 90.400 147.735 90.570 ;
        RECT 147.925 90.400 148.095 90.570 ;
        RECT 148.285 90.400 148.455 90.570 ;
        RECT 148.645 90.400 148.815 90.570 ;
        RECT 149.005 90.400 149.175 90.570 ;
        RECT 194.200 90.400 194.370 90.570 ;
        RECT 194.560 90.400 194.730 90.570 ;
        RECT 194.920 90.400 195.090 90.570 ;
        RECT 195.280 90.400 195.450 90.570 ;
        RECT 195.640 90.400 195.810 90.570 ;
        RECT 196.000 90.400 196.170 90.570 ;
        RECT 215.545 90.445 215.715 90.615 ;
        RECT 219.175 90.435 219.345 90.605 ;
        RECT 225.095 90.620 225.265 90.790 ;
        RECT 225.455 90.620 225.625 90.790 ;
        RECT 225.815 90.620 225.985 90.790 ;
        RECT 226.175 90.620 226.345 90.790 ;
        RECT 226.535 90.620 226.705 90.790 ;
        RECT 226.895 90.620 227.065 90.790 ;
        RECT 272.090 90.620 272.260 90.790 ;
        RECT 272.450 90.620 272.620 90.790 ;
        RECT 272.810 90.620 272.980 90.790 ;
        RECT 273.170 90.620 273.340 90.790 ;
        RECT 273.530 90.620 273.700 90.790 ;
        RECT 273.890 90.620 274.060 90.790 ;
        RECT 212.370 90.050 212.540 90.220 ;
        RECT 147.205 89.570 147.375 89.740 ;
        RECT 147.565 89.570 147.735 89.740 ;
        RECT 147.925 89.570 148.095 89.740 ;
        RECT 148.285 89.570 148.455 89.740 ;
        RECT 148.645 89.570 148.815 89.740 ;
        RECT 149.005 89.570 149.175 89.740 ;
        RECT 194.200 89.570 194.370 89.740 ;
        RECT 194.560 89.570 194.730 89.740 ;
        RECT 194.920 89.570 195.090 89.740 ;
        RECT 195.280 89.570 195.450 89.740 ;
        RECT 195.640 89.570 195.810 89.740 ;
        RECT 196.000 89.570 196.170 89.740 ;
        RECT 225.095 89.790 225.265 89.960 ;
        RECT 225.455 89.790 225.625 89.960 ;
        RECT 225.815 89.790 225.985 89.960 ;
        RECT 226.175 89.790 226.345 89.960 ;
        RECT 226.535 89.790 226.705 89.960 ;
        RECT 226.895 89.790 227.065 89.960 ;
        RECT 272.090 89.790 272.260 89.960 ;
        RECT 272.450 89.790 272.620 89.960 ;
        RECT 272.810 89.790 272.980 89.960 ;
        RECT 273.170 89.790 273.340 89.960 ;
        RECT 273.530 89.790 273.700 89.960 ;
        RECT 273.890 89.790 274.060 89.960 ;
        RECT 208.080 89.460 208.250 89.630 ;
        RECT 204.520 89.065 204.690 89.235 ;
        RECT 147.205 88.740 147.375 88.910 ;
        RECT 147.565 88.740 147.735 88.910 ;
        RECT 147.925 88.740 148.095 88.910 ;
        RECT 148.285 88.740 148.455 88.910 ;
        RECT 148.645 88.740 148.815 88.910 ;
        RECT 149.005 88.740 149.175 88.910 ;
        RECT 194.200 88.740 194.370 88.910 ;
        RECT 194.560 88.740 194.730 88.910 ;
        RECT 194.920 88.740 195.090 88.910 ;
        RECT 195.280 88.740 195.450 88.910 ;
        RECT 195.640 88.740 195.810 88.910 ;
        RECT 196.000 88.740 196.170 88.910 ;
        RECT 225.095 88.960 225.265 89.130 ;
        RECT 225.455 88.960 225.625 89.130 ;
        RECT 225.815 88.960 225.985 89.130 ;
        RECT 226.175 88.960 226.345 89.130 ;
        RECT 226.535 88.960 226.705 89.130 ;
        RECT 226.895 88.960 227.065 89.130 ;
        RECT 272.090 88.960 272.260 89.130 ;
        RECT 272.450 88.960 272.620 89.130 ;
        RECT 272.810 88.960 272.980 89.130 ;
        RECT 273.170 88.960 273.340 89.130 ;
        RECT 273.530 88.960 273.700 89.130 ;
        RECT 273.890 88.960 274.060 89.130 ;
        RECT 205.050 88.670 205.220 88.840 ;
        RECT 208.080 88.670 208.250 88.840 ;
        RECT 147.205 87.910 147.375 88.080 ;
        RECT 147.565 87.910 147.735 88.080 ;
        RECT 147.925 87.910 148.095 88.080 ;
        RECT 148.285 87.910 148.455 88.080 ;
        RECT 148.645 87.910 148.815 88.080 ;
        RECT 149.005 87.910 149.175 88.080 ;
        RECT 194.200 87.910 194.370 88.080 ;
        RECT 194.560 87.910 194.730 88.080 ;
        RECT 194.920 87.910 195.090 88.080 ;
        RECT 195.280 87.910 195.450 88.080 ;
        RECT 195.640 87.910 195.810 88.080 ;
        RECT 196.000 87.910 196.170 88.080 ;
        RECT 212.370 88.060 212.540 88.230 ;
        RECT 215.060 88.060 215.230 88.230 ;
        RECT 218.690 88.050 218.860 88.220 ;
        RECT 225.095 88.130 225.265 88.300 ;
        RECT 225.455 88.130 225.625 88.300 ;
        RECT 225.815 88.130 225.985 88.300 ;
        RECT 226.175 88.130 226.345 88.300 ;
        RECT 226.535 88.130 226.705 88.300 ;
        RECT 226.895 88.130 227.065 88.300 ;
        RECT 272.090 88.130 272.260 88.300 ;
        RECT 272.450 88.130 272.620 88.300 ;
        RECT 272.810 88.130 272.980 88.300 ;
        RECT 273.170 88.130 273.340 88.300 ;
        RECT 273.530 88.130 273.700 88.300 ;
        RECT 273.890 88.130 274.060 88.300 ;
        RECT 211.885 87.665 212.055 87.835 ;
        RECT 215.545 87.665 215.715 87.835 ;
        RECT 219.175 87.655 219.345 87.825 ;
        RECT 147.205 87.080 147.375 87.250 ;
        RECT 147.565 87.080 147.735 87.250 ;
        RECT 147.925 87.080 148.095 87.250 ;
        RECT 148.285 87.080 148.455 87.250 ;
        RECT 148.645 87.080 148.815 87.250 ;
        RECT 149.005 87.080 149.175 87.250 ;
        RECT 212.370 87.270 212.540 87.440 ;
        RECT 225.095 87.300 225.265 87.470 ;
        RECT 225.455 87.300 225.625 87.470 ;
        RECT 225.815 87.300 225.985 87.470 ;
        RECT 226.175 87.300 226.345 87.470 ;
        RECT 226.535 87.300 226.705 87.470 ;
        RECT 226.895 87.300 227.065 87.470 ;
        RECT 194.200 87.080 194.370 87.250 ;
        RECT 194.560 87.080 194.730 87.250 ;
        RECT 194.920 87.080 195.090 87.250 ;
        RECT 195.280 87.080 195.450 87.250 ;
        RECT 195.640 87.080 195.810 87.250 ;
        RECT 196.000 87.080 196.170 87.250 ;
        RECT 272.090 87.300 272.260 87.470 ;
        RECT 272.450 87.300 272.620 87.470 ;
        RECT 272.810 87.300 272.980 87.470 ;
        RECT 273.170 87.300 273.340 87.470 ;
        RECT 273.530 87.300 273.700 87.470 ;
        RECT 273.890 87.300 274.060 87.470 ;
        RECT 147.205 86.250 147.375 86.420 ;
        RECT 147.565 86.250 147.735 86.420 ;
        RECT 147.925 86.250 148.095 86.420 ;
        RECT 148.285 86.250 148.455 86.420 ;
        RECT 148.645 86.250 148.815 86.420 ;
        RECT 149.005 86.250 149.175 86.420 ;
        RECT 194.200 86.250 194.370 86.420 ;
        RECT 194.560 86.250 194.730 86.420 ;
        RECT 194.920 86.250 195.090 86.420 ;
        RECT 195.280 86.250 195.450 86.420 ;
        RECT 195.640 86.250 195.810 86.420 ;
        RECT 196.000 86.250 196.170 86.420 ;
        RECT 205.050 86.380 205.220 86.550 ;
        RECT 208.080 86.380 208.250 86.550 ;
        RECT 225.095 86.470 225.265 86.640 ;
        RECT 225.455 86.470 225.625 86.640 ;
        RECT 225.815 86.470 225.985 86.640 ;
        RECT 226.175 86.470 226.345 86.640 ;
        RECT 226.535 86.470 226.705 86.640 ;
        RECT 226.895 86.470 227.065 86.640 ;
        RECT 272.090 86.470 272.260 86.640 ;
        RECT 272.450 86.470 272.620 86.640 ;
        RECT 272.810 86.470 272.980 86.640 ;
        RECT 273.170 86.470 273.340 86.640 ;
        RECT 273.530 86.470 273.700 86.640 ;
        RECT 273.890 86.470 274.060 86.640 ;
        RECT 204.520 85.985 204.690 86.155 ;
        RECT 208.610 85.985 208.780 86.155 ;
        RECT 147.205 85.420 147.375 85.590 ;
        RECT 147.565 85.420 147.735 85.590 ;
        RECT 147.925 85.420 148.095 85.590 ;
        RECT 148.285 85.420 148.455 85.590 ;
        RECT 148.645 85.420 148.815 85.590 ;
        RECT 149.005 85.420 149.175 85.590 ;
        RECT 194.200 85.420 194.370 85.590 ;
        RECT 194.560 85.420 194.730 85.590 ;
        RECT 194.920 85.420 195.090 85.590 ;
        RECT 195.280 85.420 195.450 85.590 ;
        RECT 195.640 85.420 195.810 85.590 ;
        RECT 196.000 85.420 196.170 85.590 ;
        RECT 225.095 85.640 225.265 85.810 ;
        RECT 225.455 85.640 225.625 85.810 ;
        RECT 225.815 85.640 225.985 85.810 ;
        RECT 226.175 85.640 226.345 85.810 ;
        RECT 226.535 85.640 226.705 85.810 ;
        RECT 226.895 85.640 227.065 85.810 ;
        RECT 272.090 85.640 272.260 85.810 ;
        RECT 272.450 85.640 272.620 85.810 ;
        RECT 272.810 85.640 272.980 85.810 ;
        RECT 273.170 85.640 273.340 85.810 ;
        RECT 273.530 85.640 273.700 85.810 ;
        RECT 273.890 85.640 274.060 85.810 ;
        RECT 212.370 85.280 212.540 85.450 ;
        RECT 215.060 85.280 215.230 85.450 ;
        RECT 218.690 85.270 218.860 85.440 ;
        RECT 211.885 84.885 212.055 85.055 ;
        RECT 194.200 84.590 194.370 84.760 ;
        RECT 194.560 84.590 194.730 84.760 ;
        RECT 194.920 84.590 195.090 84.760 ;
        RECT 195.280 84.590 195.450 84.760 ;
        RECT 195.640 84.590 195.810 84.760 ;
        RECT 196.000 84.590 196.170 84.760 ;
        RECT 215.545 84.885 215.715 85.055 ;
        RECT 219.175 84.875 219.345 85.045 ;
        RECT 225.095 84.810 225.265 84.980 ;
        RECT 225.455 84.810 225.625 84.980 ;
        RECT 225.815 84.810 225.985 84.980 ;
        RECT 226.175 84.810 226.345 84.980 ;
        RECT 226.535 84.810 226.705 84.980 ;
        RECT 226.895 84.810 227.065 84.980 ;
        RECT 272.090 84.810 272.260 84.980 ;
        RECT 272.450 84.810 272.620 84.980 ;
        RECT 272.810 84.810 272.980 84.980 ;
        RECT 273.170 84.810 273.340 84.980 ;
        RECT 273.530 84.810 273.700 84.980 ;
        RECT 273.890 84.810 274.060 84.980 ;
        RECT 212.370 84.490 212.540 84.660 ;
        RECT 218.690 84.480 218.860 84.650 ;
        RECT 225.095 83.980 225.265 84.150 ;
        RECT 225.455 83.980 225.625 84.150 ;
        RECT 225.815 83.980 225.985 84.150 ;
        RECT 226.175 83.980 226.345 84.150 ;
        RECT 226.535 83.980 226.705 84.150 ;
        RECT 226.895 83.980 227.065 84.150 ;
        RECT 272.090 83.980 272.260 84.150 ;
        RECT 272.450 83.980 272.620 84.150 ;
        RECT 272.810 83.980 272.980 84.150 ;
        RECT 273.170 83.980 273.340 84.150 ;
        RECT 273.530 83.980 273.700 84.150 ;
        RECT 273.890 83.980 274.060 84.150 ;
        RECT 225.095 83.150 225.265 83.320 ;
        RECT 225.455 83.150 225.625 83.320 ;
        RECT 225.815 83.150 225.985 83.320 ;
        RECT 226.175 83.150 226.345 83.320 ;
        RECT 226.535 83.150 226.705 83.320 ;
        RECT 226.895 83.150 227.065 83.320 ;
        RECT 272.090 83.150 272.260 83.320 ;
        RECT 272.450 83.150 272.620 83.320 ;
        RECT 272.810 83.150 272.980 83.320 ;
        RECT 273.170 83.150 273.340 83.320 ;
        RECT 273.530 83.150 273.700 83.320 ;
        RECT 273.890 83.150 274.060 83.320 ;
        RECT 225.095 82.320 225.265 82.490 ;
        RECT 225.455 82.320 225.625 82.490 ;
        RECT 225.815 82.320 225.985 82.490 ;
        RECT 226.175 82.320 226.345 82.490 ;
        RECT 226.535 82.320 226.705 82.490 ;
        RECT 226.895 82.320 227.065 82.490 ;
        RECT 272.090 82.320 272.260 82.490 ;
        RECT 272.450 82.320 272.620 82.490 ;
        RECT 272.810 82.320 272.980 82.490 ;
        RECT 273.170 82.320 273.340 82.490 ;
        RECT 273.530 82.320 273.700 82.490 ;
        RECT 273.890 82.320 274.060 82.490 ;
        RECT 147.255 81.590 147.425 81.760 ;
        RECT 147.615 81.590 147.785 81.760 ;
        RECT 147.975 81.590 148.145 81.760 ;
        RECT 148.335 81.590 148.505 81.760 ;
        RECT 148.695 81.590 148.865 81.760 ;
        RECT 149.055 81.590 149.225 81.760 ;
        RECT 194.250 81.590 194.420 81.760 ;
        RECT 194.610 81.590 194.780 81.760 ;
        RECT 194.970 81.590 195.140 81.760 ;
        RECT 195.330 81.590 195.500 81.760 ;
        RECT 195.690 81.590 195.860 81.760 ;
        RECT 196.050 81.590 196.220 81.760 ;
        RECT 225.095 81.490 225.265 81.660 ;
        RECT 225.455 81.490 225.625 81.660 ;
        RECT 225.815 81.490 225.985 81.660 ;
        RECT 226.175 81.490 226.345 81.660 ;
        RECT 226.535 81.490 226.705 81.660 ;
        RECT 226.895 81.490 227.065 81.660 ;
        RECT 272.090 81.490 272.260 81.660 ;
        RECT 272.450 81.490 272.620 81.660 ;
        RECT 272.810 81.490 272.980 81.660 ;
        RECT 273.170 81.490 273.340 81.660 ;
        RECT 273.530 81.490 273.700 81.660 ;
        RECT 273.890 81.490 274.060 81.660 ;
        RECT 147.255 80.760 147.425 80.930 ;
        RECT 147.615 80.760 147.785 80.930 ;
        RECT 147.975 80.760 148.145 80.930 ;
        RECT 148.335 80.760 148.505 80.930 ;
        RECT 148.695 80.760 148.865 80.930 ;
        RECT 149.055 80.760 149.225 80.930 ;
        RECT 194.250 80.760 194.420 80.930 ;
        RECT 194.610 80.760 194.780 80.930 ;
        RECT 194.970 80.760 195.140 80.930 ;
        RECT 195.330 80.760 195.500 80.930 ;
        RECT 195.690 80.760 195.860 80.930 ;
        RECT 196.050 80.760 196.220 80.930 ;
        RECT 225.095 80.660 225.265 80.830 ;
        RECT 225.455 80.660 225.625 80.830 ;
        RECT 225.815 80.660 225.985 80.830 ;
        RECT 226.175 80.660 226.345 80.830 ;
        RECT 226.535 80.660 226.705 80.830 ;
        RECT 226.895 80.660 227.065 80.830 ;
        RECT 272.090 80.660 272.260 80.830 ;
        RECT 272.450 80.660 272.620 80.830 ;
        RECT 272.810 80.660 272.980 80.830 ;
        RECT 273.170 80.660 273.340 80.830 ;
        RECT 273.530 80.660 273.700 80.830 ;
        RECT 273.890 80.660 274.060 80.830 ;
        RECT 147.255 79.930 147.425 80.100 ;
        RECT 147.615 79.930 147.785 80.100 ;
        RECT 147.975 79.930 148.145 80.100 ;
        RECT 148.335 79.930 148.505 80.100 ;
        RECT 148.695 79.930 148.865 80.100 ;
        RECT 149.055 79.930 149.225 80.100 ;
        RECT 194.250 79.930 194.420 80.100 ;
        RECT 194.610 79.930 194.780 80.100 ;
        RECT 194.970 79.930 195.140 80.100 ;
        RECT 195.330 79.930 195.500 80.100 ;
        RECT 195.690 79.930 195.860 80.100 ;
        RECT 196.050 79.930 196.220 80.100 ;
        RECT 147.255 79.100 147.425 79.270 ;
        RECT 147.615 79.100 147.785 79.270 ;
        RECT 147.975 79.100 148.145 79.270 ;
        RECT 148.335 79.100 148.505 79.270 ;
        RECT 148.695 79.100 148.865 79.270 ;
        RECT 149.055 79.100 149.225 79.270 ;
        RECT 194.250 79.100 194.420 79.270 ;
        RECT 194.610 79.100 194.780 79.270 ;
        RECT 194.970 79.100 195.140 79.270 ;
        RECT 195.330 79.100 195.500 79.270 ;
        RECT 195.690 79.100 195.860 79.270 ;
        RECT 196.050 79.100 196.220 79.270 ;
        RECT 147.255 78.270 147.425 78.440 ;
        RECT 147.615 78.270 147.785 78.440 ;
        RECT 147.975 78.270 148.145 78.440 ;
        RECT 148.335 78.270 148.505 78.440 ;
        RECT 148.695 78.270 148.865 78.440 ;
        RECT 149.055 78.270 149.225 78.440 ;
        RECT 194.250 78.270 194.420 78.440 ;
        RECT 194.610 78.270 194.780 78.440 ;
        RECT 194.970 78.270 195.140 78.440 ;
        RECT 195.330 78.270 195.500 78.440 ;
        RECT 195.690 78.270 195.860 78.440 ;
        RECT 196.050 78.270 196.220 78.440 ;
        RECT 147.255 77.440 147.425 77.610 ;
        RECT 147.615 77.440 147.785 77.610 ;
        RECT 147.975 77.440 148.145 77.610 ;
        RECT 148.335 77.440 148.505 77.610 ;
        RECT 148.695 77.440 148.865 77.610 ;
        RECT 149.055 77.440 149.225 77.610 ;
        RECT 194.250 77.440 194.420 77.610 ;
        RECT 194.610 77.440 194.780 77.610 ;
        RECT 194.970 77.440 195.140 77.610 ;
        RECT 195.330 77.440 195.500 77.610 ;
        RECT 195.690 77.440 195.860 77.610 ;
        RECT 196.050 77.440 196.220 77.610 ;
        RECT 147.255 76.610 147.425 76.780 ;
        RECT 147.615 76.610 147.785 76.780 ;
        RECT 147.975 76.610 148.145 76.780 ;
        RECT 148.335 76.610 148.505 76.780 ;
        RECT 148.695 76.610 148.865 76.780 ;
        RECT 149.055 76.610 149.225 76.780 ;
        RECT 194.250 76.610 194.420 76.780 ;
        RECT 194.610 76.610 194.780 76.780 ;
        RECT 194.970 76.610 195.140 76.780 ;
        RECT 195.330 76.610 195.500 76.780 ;
        RECT 195.690 76.610 195.860 76.780 ;
        RECT 196.050 76.610 196.220 76.780 ;
        RECT 147.255 75.780 147.425 75.950 ;
        RECT 147.615 75.780 147.785 75.950 ;
        RECT 147.975 75.780 148.145 75.950 ;
        RECT 148.335 75.780 148.505 75.950 ;
        RECT 148.695 75.780 148.865 75.950 ;
        RECT 149.055 75.780 149.225 75.950 ;
        RECT 194.250 75.780 194.420 75.950 ;
        RECT 194.610 75.780 194.780 75.950 ;
        RECT 194.970 75.780 195.140 75.950 ;
        RECT 195.330 75.780 195.500 75.950 ;
        RECT 195.690 75.780 195.860 75.950 ;
        RECT 196.050 75.780 196.220 75.950 ;
        RECT 147.255 74.950 147.425 75.120 ;
        RECT 147.615 74.950 147.785 75.120 ;
        RECT 147.975 74.950 148.145 75.120 ;
        RECT 148.335 74.950 148.505 75.120 ;
        RECT 148.695 74.950 148.865 75.120 ;
        RECT 149.055 74.950 149.225 75.120 ;
        RECT 194.250 74.950 194.420 75.120 ;
        RECT 194.610 74.950 194.780 75.120 ;
        RECT 194.970 74.950 195.140 75.120 ;
        RECT 195.330 74.950 195.500 75.120 ;
        RECT 195.690 74.950 195.860 75.120 ;
        RECT 196.050 74.950 196.220 75.120 ;
        RECT 205.100 79.100 205.270 79.270 ;
        RECT 208.450 79.100 208.620 79.270 ;
        RECT 212.960 79.100 213.130 79.270 ;
        RECT 216.310 79.100 216.480 79.270 ;
        RECT 201.120 78.695 201.290 78.865 ;
        RECT 202.090 78.695 202.260 78.865 ;
        RECT 204.570 78.705 204.740 78.875 ;
        RECT 205.630 78.705 205.800 78.875 ;
        RECT 207.920 78.705 208.090 78.875 ;
        RECT 208.980 78.705 209.150 78.875 ;
        RECT 212.430 78.705 212.600 78.875 ;
        RECT 213.490 78.705 213.660 78.875 ;
        RECT 215.780 78.705 215.950 78.875 ;
        RECT 216.840 78.705 217.010 78.875 ;
        RECT 219.320 78.695 219.490 78.865 ;
        RECT 220.290 78.695 220.460 78.865 ;
        RECT 201.605 78.300 201.775 78.470 ;
        RECT 205.100 78.310 205.270 78.480 ;
        RECT 216.310 78.310 216.480 78.480 ;
        RECT 219.805 78.300 219.975 78.470 ;
        RECT 201.595 76.060 201.765 76.230 ;
        RECT 205.110 76.050 205.280 76.220 ;
        RECT 216.300 76.050 216.470 76.220 ;
        RECT 219.815 76.060 219.985 76.230 ;
        RECT 204.580 75.655 204.750 75.825 ;
        RECT 205.640 75.655 205.810 75.825 ;
        RECT 207.920 75.625 208.090 75.795 ;
        RECT 208.980 75.625 209.150 75.795 ;
        RECT 212.430 75.625 212.600 75.795 ;
        RECT 213.490 75.625 213.660 75.795 ;
        RECT 215.770 75.655 215.940 75.825 ;
        RECT 216.830 75.655 217.000 75.825 ;
        RECT 205.110 75.260 205.280 75.430 ;
        RECT 208.450 75.230 208.620 75.400 ;
        RECT 212.960 75.230 213.130 75.400 ;
        RECT 216.300 75.260 216.470 75.430 ;
        RECT 225.095 79.830 225.265 80.000 ;
        RECT 225.455 79.830 225.625 80.000 ;
        RECT 225.815 79.830 225.985 80.000 ;
        RECT 226.175 79.830 226.345 80.000 ;
        RECT 226.535 79.830 226.705 80.000 ;
        RECT 226.895 79.830 227.065 80.000 ;
        RECT 272.090 79.830 272.260 80.000 ;
        RECT 272.450 79.830 272.620 80.000 ;
        RECT 272.810 79.830 272.980 80.000 ;
        RECT 273.170 79.830 273.340 80.000 ;
        RECT 273.530 79.830 273.700 80.000 ;
        RECT 273.890 79.830 274.060 80.000 ;
        RECT 225.095 79.000 225.265 79.170 ;
        RECT 225.455 79.000 225.625 79.170 ;
        RECT 225.815 79.000 225.985 79.170 ;
        RECT 226.175 79.000 226.345 79.170 ;
        RECT 226.535 79.000 226.705 79.170 ;
        RECT 226.895 79.000 227.065 79.170 ;
        RECT 272.090 79.000 272.260 79.170 ;
        RECT 272.450 79.000 272.620 79.170 ;
        RECT 272.810 79.000 272.980 79.170 ;
        RECT 273.170 79.000 273.340 79.170 ;
        RECT 273.530 79.000 273.700 79.170 ;
        RECT 273.890 79.000 274.060 79.170 ;
        RECT 225.095 78.170 225.265 78.340 ;
        RECT 225.455 78.170 225.625 78.340 ;
        RECT 225.815 78.170 225.985 78.340 ;
        RECT 226.175 78.170 226.345 78.340 ;
        RECT 226.535 78.170 226.705 78.340 ;
        RECT 226.895 78.170 227.065 78.340 ;
        RECT 272.090 78.170 272.260 78.340 ;
        RECT 272.450 78.170 272.620 78.340 ;
        RECT 272.810 78.170 272.980 78.340 ;
        RECT 273.170 78.170 273.340 78.340 ;
        RECT 273.530 78.170 273.700 78.340 ;
        RECT 273.890 78.170 274.060 78.340 ;
        RECT 225.095 77.340 225.265 77.510 ;
        RECT 225.455 77.340 225.625 77.510 ;
        RECT 225.815 77.340 225.985 77.510 ;
        RECT 226.175 77.340 226.345 77.510 ;
        RECT 226.535 77.340 226.705 77.510 ;
        RECT 226.895 77.340 227.065 77.510 ;
        RECT 272.090 77.340 272.260 77.510 ;
        RECT 272.450 77.340 272.620 77.510 ;
        RECT 272.810 77.340 272.980 77.510 ;
        RECT 273.170 77.340 273.340 77.510 ;
        RECT 273.530 77.340 273.700 77.510 ;
        RECT 273.890 77.340 274.060 77.510 ;
        RECT 225.095 76.510 225.265 76.680 ;
        RECT 225.455 76.510 225.625 76.680 ;
        RECT 225.815 76.510 225.985 76.680 ;
        RECT 226.175 76.510 226.345 76.680 ;
        RECT 226.535 76.510 226.705 76.680 ;
        RECT 226.895 76.510 227.065 76.680 ;
        RECT 272.090 76.510 272.260 76.680 ;
        RECT 272.450 76.510 272.620 76.680 ;
        RECT 272.810 76.510 272.980 76.680 ;
        RECT 273.170 76.510 273.340 76.680 ;
        RECT 273.530 76.510 273.700 76.680 ;
        RECT 273.890 76.510 274.060 76.680 ;
        RECT 225.095 75.680 225.265 75.850 ;
        RECT 225.455 75.680 225.625 75.850 ;
        RECT 225.815 75.680 225.985 75.850 ;
        RECT 226.175 75.680 226.345 75.850 ;
        RECT 226.535 75.680 226.705 75.850 ;
        RECT 226.895 75.680 227.065 75.850 ;
        RECT 272.090 75.680 272.260 75.850 ;
        RECT 272.450 75.680 272.620 75.850 ;
        RECT 272.810 75.680 272.980 75.850 ;
        RECT 273.170 75.680 273.340 75.850 ;
        RECT 273.530 75.680 273.700 75.850 ;
        RECT 273.890 75.680 274.060 75.850 ;
        RECT 225.095 74.850 225.265 75.020 ;
        RECT 225.455 74.850 225.625 75.020 ;
        RECT 225.815 74.850 225.985 75.020 ;
        RECT 226.175 74.850 226.345 75.020 ;
        RECT 226.535 74.850 226.705 75.020 ;
        RECT 226.895 74.850 227.065 75.020 ;
        RECT 272.090 74.850 272.260 75.020 ;
        RECT 272.450 74.850 272.620 75.020 ;
        RECT 272.810 74.850 272.980 75.020 ;
        RECT 273.170 74.850 273.340 75.020 ;
        RECT 273.530 74.850 273.700 75.020 ;
        RECT 273.890 74.850 274.060 75.020 ;
        RECT 147.255 74.120 147.425 74.290 ;
        RECT 147.615 74.120 147.785 74.290 ;
        RECT 147.975 74.120 148.145 74.290 ;
        RECT 148.335 74.120 148.505 74.290 ;
        RECT 148.695 74.120 148.865 74.290 ;
        RECT 149.055 74.120 149.225 74.290 ;
        RECT 194.250 74.120 194.420 74.290 ;
        RECT 194.610 74.120 194.780 74.290 ;
        RECT 194.970 74.120 195.140 74.290 ;
        RECT 195.330 74.120 195.500 74.290 ;
        RECT 195.690 74.120 195.860 74.290 ;
        RECT 196.050 74.120 196.220 74.290 ;
        RECT 225.095 74.020 225.265 74.190 ;
        RECT 225.455 74.020 225.625 74.190 ;
        RECT 225.815 74.020 225.985 74.190 ;
        RECT 226.175 74.020 226.345 74.190 ;
        RECT 226.535 74.020 226.705 74.190 ;
        RECT 226.895 74.020 227.065 74.190 ;
        RECT 272.090 74.020 272.260 74.190 ;
        RECT 272.450 74.020 272.620 74.190 ;
        RECT 272.810 74.020 272.980 74.190 ;
        RECT 273.170 74.020 273.340 74.190 ;
        RECT 273.530 74.020 273.700 74.190 ;
        RECT 273.890 74.020 274.060 74.190 ;
        RECT 147.255 73.290 147.425 73.460 ;
        RECT 147.615 73.290 147.785 73.460 ;
        RECT 147.975 73.290 148.145 73.460 ;
        RECT 148.335 73.290 148.505 73.460 ;
        RECT 148.695 73.290 148.865 73.460 ;
        RECT 149.055 73.290 149.225 73.460 ;
        RECT 194.250 73.290 194.420 73.460 ;
        RECT 194.610 73.290 194.780 73.460 ;
        RECT 194.970 73.290 195.140 73.460 ;
        RECT 195.330 73.290 195.500 73.460 ;
        RECT 195.690 73.290 195.860 73.460 ;
        RECT 196.050 73.290 196.220 73.460 ;
        RECT 225.095 73.190 225.265 73.360 ;
        RECT 225.455 73.190 225.625 73.360 ;
        RECT 225.815 73.190 225.985 73.360 ;
        RECT 226.175 73.190 226.345 73.360 ;
        RECT 226.535 73.190 226.705 73.360 ;
        RECT 226.895 73.190 227.065 73.360 ;
        RECT 272.090 73.190 272.260 73.360 ;
        RECT 272.450 73.190 272.620 73.360 ;
        RECT 272.810 73.190 272.980 73.360 ;
        RECT 273.170 73.190 273.340 73.360 ;
        RECT 273.530 73.190 273.700 73.360 ;
        RECT 273.890 73.190 274.060 73.360 ;
        RECT 147.255 72.460 147.425 72.630 ;
        RECT 147.615 72.460 147.785 72.630 ;
        RECT 147.975 72.460 148.145 72.630 ;
        RECT 148.335 72.460 148.505 72.630 ;
        RECT 148.695 72.460 148.865 72.630 ;
        RECT 149.055 72.460 149.225 72.630 ;
        RECT 194.250 72.460 194.420 72.630 ;
        RECT 194.610 72.460 194.780 72.630 ;
        RECT 194.970 72.460 195.140 72.630 ;
        RECT 195.330 72.460 195.500 72.630 ;
        RECT 195.690 72.460 195.860 72.630 ;
        RECT 196.050 72.460 196.220 72.630 ;
        RECT 225.095 72.360 225.265 72.530 ;
        RECT 225.455 72.360 225.625 72.530 ;
        RECT 225.815 72.360 225.985 72.530 ;
        RECT 226.175 72.360 226.345 72.530 ;
        RECT 226.535 72.360 226.705 72.530 ;
        RECT 226.895 72.360 227.065 72.530 ;
        RECT 272.090 72.360 272.260 72.530 ;
        RECT 272.450 72.360 272.620 72.530 ;
        RECT 272.810 72.360 272.980 72.530 ;
        RECT 273.170 72.360 273.340 72.530 ;
        RECT 273.530 72.360 273.700 72.530 ;
        RECT 273.890 72.360 274.060 72.530 ;
        RECT 147.255 71.630 147.425 71.800 ;
        RECT 147.615 71.630 147.785 71.800 ;
        RECT 147.975 71.630 148.145 71.800 ;
        RECT 148.335 71.630 148.505 71.800 ;
        RECT 148.695 71.630 148.865 71.800 ;
        RECT 149.055 71.630 149.225 71.800 ;
        RECT 194.250 71.630 194.420 71.800 ;
        RECT 194.610 71.630 194.780 71.800 ;
        RECT 194.970 71.630 195.140 71.800 ;
        RECT 195.330 71.630 195.500 71.800 ;
        RECT 195.690 71.630 195.860 71.800 ;
        RECT 196.050 71.630 196.220 71.800 ;
        RECT 225.095 71.530 225.265 71.700 ;
        RECT 225.455 71.530 225.625 71.700 ;
        RECT 225.815 71.530 225.985 71.700 ;
        RECT 226.175 71.530 226.345 71.700 ;
        RECT 226.535 71.530 226.705 71.700 ;
        RECT 226.895 71.530 227.065 71.700 ;
        RECT 272.090 71.530 272.260 71.700 ;
        RECT 272.450 71.530 272.620 71.700 ;
        RECT 272.810 71.530 272.980 71.700 ;
        RECT 273.170 71.530 273.340 71.700 ;
        RECT 273.530 71.530 273.700 71.700 ;
        RECT 273.890 71.530 274.060 71.700 ;
        RECT 147.255 70.800 147.425 70.970 ;
        RECT 147.615 70.800 147.785 70.970 ;
        RECT 147.975 70.800 148.145 70.970 ;
        RECT 148.335 70.800 148.505 70.970 ;
        RECT 148.695 70.800 148.865 70.970 ;
        RECT 149.055 70.800 149.225 70.970 ;
        RECT 194.250 70.800 194.420 70.970 ;
        RECT 194.610 70.800 194.780 70.970 ;
        RECT 194.970 70.800 195.140 70.970 ;
        RECT 195.330 70.800 195.500 70.970 ;
        RECT 195.690 70.800 195.860 70.970 ;
        RECT 196.050 70.800 196.220 70.970 ;
        RECT 215.885 70.400 217.855 70.930 ;
        RECT 225.095 70.700 225.265 70.870 ;
        RECT 225.455 70.700 225.625 70.870 ;
        RECT 225.815 70.700 225.985 70.870 ;
        RECT 226.175 70.700 226.345 70.870 ;
        RECT 226.535 70.700 226.705 70.870 ;
        RECT 226.895 70.700 227.065 70.870 ;
        RECT 272.090 70.700 272.260 70.870 ;
        RECT 272.450 70.700 272.620 70.870 ;
        RECT 272.810 70.700 272.980 70.870 ;
        RECT 273.170 70.700 273.340 70.870 ;
        RECT 273.530 70.700 273.700 70.870 ;
        RECT 273.890 70.700 274.060 70.870 ;
        RECT 147.255 69.970 147.425 70.140 ;
        RECT 147.615 69.970 147.785 70.140 ;
        RECT 147.975 69.970 148.145 70.140 ;
        RECT 148.335 69.970 148.505 70.140 ;
        RECT 148.695 69.970 148.865 70.140 ;
        RECT 149.055 69.970 149.225 70.140 ;
        RECT 194.250 69.970 194.420 70.140 ;
        RECT 194.610 69.970 194.780 70.140 ;
        RECT 194.970 69.970 195.140 70.140 ;
        RECT 195.330 69.970 195.500 70.140 ;
        RECT 195.690 69.970 195.860 70.140 ;
        RECT 196.050 69.970 196.220 70.140 ;
        RECT 225.095 69.870 225.265 70.040 ;
        RECT 225.455 69.870 225.625 70.040 ;
        RECT 225.815 69.870 225.985 70.040 ;
        RECT 226.175 69.870 226.345 70.040 ;
        RECT 226.535 69.870 226.705 70.040 ;
        RECT 226.895 69.870 227.065 70.040 ;
        RECT 272.090 69.870 272.260 70.040 ;
        RECT 272.450 69.870 272.620 70.040 ;
        RECT 272.810 69.870 272.980 70.040 ;
        RECT 273.170 69.870 273.340 70.040 ;
        RECT 273.530 69.870 273.700 70.040 ;
        RECT 273.890 69.870 274.060 70.040 ;
        RECT 147.255 69.140 147.425 69.310 ;
        RECT 147.615 69.140 147.785 69.310 ;
        RECT 147.975 69.140 148.145 69.310 ;
        RECT 148.335 69.140 148.505 69.310 ;
        RECT 148.695 69.140 148.865 69.310 ;
        RECT 149.055 69.140 149.225 69.310 ;
        RECT 194.250 69.140 194.420 69.310 ;
        RECT 194.610 69.140 194.780 69.310 ;
        RECT 194.970 69.140 195.140 69.310 ;
        RECT 195.330 69.140 195.500 69.310 ;
        RECT 195.690 69.140 195.860 69.310 ;
        RECT 196.050 69.140 196.220 69.310 ;
        RECT 225.095 69.040 225.265 69.210 ;
        RECT 225.455 69.040 225.625 69.210 ;
        RECT 225.815 69.040 225.985 69.210 ;
        RECT 226.175 69.040 226.345 69.210 ;
        RECT 226.535 69.040 226.705 69.210 ;
        RECT 226.895 69.040 227.065 69.210 ;
        RECT 272.090 69.040 272.260 69.210 ;
        RECT 272.450 69.040 272.620 69.210 ;
        RECT 272.810 69.040 272.980 69.210 ;
        RECT 273.170 69.040 273.340 69.210 ;
        RECT 273.530 69.040 273.700 69.210 ;
        RECT 273.890 69.040 274.060 69.210 ;
        RECT 147.255 68.310 147.425 68.480 ;
        RECT 147.615 68.310 147.785 68.480 ;
        RECT 147.975 68.310 148.145 68.480 ;
        RECT 148.335 68.310 148.505 68.480 ;
        RECT 148.695 68.310 148.865 68.480 ;
        RECT 149.055 68.310 149.225 68.480 ;
        RECT 194.250 68.310 194.420 68.480 ;
        RECT 194.610 68.310 194.780 68.480 ;
        RECT 194.970 68.310 195.140 68.480 ;
        RECT 195.330 68.310 195.500 68.480 ;
        RECT 195.690 68.310 195.860 68.480 ;
        RECT 196.050 68.310 196.220 68.480 ;
        RECT 225.095 68.210 225.265 68.380 ;
        RECT 225.455 68.210 225.625 68.380 ;
        RECT 225.815 68.210 225.985 68.380 ;
        RECT 226.175 68.210 226.345 68.380 ;
        RECT 226.535 68.210 226.705 68.380 ;
        RECT 226.895 68.210 227.065 68.380 ;
        RECT 272.090 68.210 272.260 68.380 ;
        RECT 272.450 68.210 272.620 68.380 ;
        RECT 272.810 68.210 272.980 68.380 ;
        RECT 273.170 68.210 273.340 68.380 ;
        RECT 273.530 68.210 273.700 68.380 ;
        RECT 273.890 68.210 274.060 68.380 ;
        RECT 147.255 67.480 147.425 67.650 ;
        RECT 147.615 67.480 147.785 67.650 ;
        RECT 147.975 67.480 148.145 67.650 ;
        RECT 148.335 67.480 148.505 67.650 ;
        RECT 148.695 67.480 148.865 67.650 ;
        RECT 149.055 67.480 149.225 67.650 ;
        RECT 194.250 67.480 194.420 67.650 ;
        RECT 194.610 67.480 194.780 67.650 ;
        RECT 194.970 67.480 195.140 67.650 ;
        RECT 195.330 67.480 195.500 67.650 ;
        RECT 195.690 67.480 195.860 67.650 ;
        RECT 196.050 67.480 196.220 67.650 ;
        RECT 203.035 67.610 203.205 67.780 ;
        RECT 203.395 67.610 203.565 67.780 ;
        RECT 206.225 67.610 206.395 67.780 ;
        RECT 206.585 67.610 206.755 67.780 ;
        RECT 214.825 67.610 214.995 67.780 ;
        RECT 215.185 67.610 215.355 67.780 ;
        RECT 218.015 67.610 218.185 67.780 ;
        RECT 218.375 67.610 218.545 67.780 ;
        RECT 225.095 67.380 225.265 67.550 ;
        RECT 225.455 67.380 225.625 67.550 ;
        RECT 225.815 67.380 225.985 67.550 ;
        RECT 226.175 67.380 226.345 67.550 ;
        RECT 226.535 67.380 226.705 67.550 ;
        RECT 226.895 67.380 227.065 67.550 ;
        RECT 272.090 67.380 272.260 67.550 ;
        RECT 272.450 67.380 272.620 67.550 ;
        RECT 272.810 67.380 272.980 67.550 ;
        RECT 273.170 67.380 273.340 67.550 ;
        RECT 273.530 67.380 273.700 67.550 ;
        RECT 273.890 67.380 274.060 67.550 ;
        RECT 209.655 66.965 209.825 67.135 ;
        RECT 194.250 66.650 194.420 66.820 ;
        RECT 194.610 66.650 194.780 66.820 ;
        RECT 194.970 66.650 195.140 66.820 ;
        RECT 195.330 66.650 195.500 66.820 ;
        RECT 195.690 66.650 195.860 66.820 ;
        RECT 196.050 66.650 196.220 66.820 ;
        RECT 210.180 66.745 210.350 66.915 ;
        RECT 225.095 66.550 225.265 66.720 ;
        RECT 225.455 66.550 225.625 66.720 ;
        RECT 225.815 66.550 225.985 66.720 ;
        RECT 226.175 66.550 226.345 66.720 ;
        RECT 226.535 66.550 226.705 66.720 ;
        RECT 226.895 66.550 227.065 66.720 ;
        RECT 272.090 66.550 272.260 66.720 ;
        RECT 272.450 66.550 272.620 66.720 ;
        RECT 272.810 66.550 272.980 66.720 ;
        RECT 273.170 66.550 273.340 66.720 ;
        RECT 273.530 66.550 273.700 66.720 ;
        RECT 273.890 66.550 274.060 66.720 ;
        RECT 210.180 65.120 210.350 65.290 ;
        RECT 206.910 64.900 207.080 65.070 ;
        RECT 205.910 64.680 206.080 64.850 ;
        RECT 206.270 64.680 206.440 64.850 ;
        RECT 211.945 64.900 212.115 65.070 ;
        RECT 210.180 64.680 210.350 64.850 ;
        RECT 212.430 64.680 212.600 64.850 ;
      LAYER met1 ;
        RECT 147.105 130.150 149.265 131.330 ;
        RECT 194.105 130.980 197.935 131.330 ;
        RECT 147.105 128.490 149.265 129.670 ;
        RECT 194.105 129.320 196.265 130.500 ;
        RECT 147.105 126.830 149.265 128.010 ;
        RECT 194.105 127.660 196.265 128.840 ;
        RECT 147.105 125.170 149.265 126.350 ;
        RECT 194.105 126.000 196.265 127.180 ;
        RECT 147.105 123.510 149.265 124.690 ;
        RECT 194.105 124.340 196.265 125.520 ;
        RECT 147.105 121.850 149.265 123.030 ;
        RECT 194.105 122.680 196.265 123.860 ;
        RECT 147.105 120.190 149.265 121.370 ;
        RECT 194.105 121.020 196.265 122.200 ;
        RECT 147.105 118.530 149.265 119.710 ;
        RECT 194.105 119.360 196.265 120.540 ;
        RECT 147.105 116.870 149.265 118.050 ;
        RECT 194.105 117.700 196.265 118.880 ;
        RECT 147.105 115.210 149.265 116.390 ;
        RECT 194.105 116.040 196.265 117.220 ;
        RECT 147.105 113.550 149.265 114.730 ;
        RECT 194.105 114.380 196.265 115.560 ;
        RECT 147.105 111.890 149.265 113.070 ;
        RECT 194.105 112.720 196.265 113.900 ;
        RECT 147.105 110.230 149.265 111.410 ;
        RECT 194.105 111.060 196.265 112.240 ;
        RECT 147.105 108.570 149.265 109.750 ;
        RECT 194.105 109.400 196.265 110.580 ;
        RECT 147.105 106.910 149.265 108.090 ;
        RECT 194.105 107.740 196.265 108.920 ;
        RECT 147.105 105.250 149.265 106.430 ;
        RECT 194.105 106.080 196.265 107.260 ;
        RECT 147.105 103.590 149.265 104.770 ;
        RECT 194.105 104.420 196.265 105.600 ;
        RECT 147.105 101.930 149.265 103.110 ;
        RECT 194.105 102.760 196.265 103.940 ;
        RECT 147.105 100.270 149.265 101.450 ;
        RECT 194.105 101.100 196.265 102.280 ;
        RECT 197.440 102.165 197.935 130.980 ;
        RECT 199.165 128.890 201.325 130.750 ;
        RECT 224.995 130.365 227.155 131.550 ;
        RECT 199.165 126.550 201.325 128.410 ;
        RECT 220.165 127.720 222.325 129.580 ;
        RECT 224.995 128.710 227.155 129.895 ;
        RECT 271.995 129.540 274.155 130.720 ;
        RECT 199.165 124.210 201.325 126.070 ;
        RECT 220.165 125.380 222.325 127.240 ;
        RECT 224.995 127.055 227.155 128.240 ;
        RECT 271.995 127.880 274.155 129.060 ;
        RECT 224.995 125.400 227.155 126.585 ;
        RECT 271.995 126.220 274.155 127.400 ;
        RECT 199.165 121.870 201.325 123.730 ;
        RECT 220.165 123.040 222.325 124.900 ;
        RECT 224.995 123.745 227.155 124.930 ;
        RECT 271.995 124.560 274.155 125.740 ;
        RECT 199.165 119.530 201.325 121.390 ;
        RECT 220.165 120.700 222.325 122.560 ;
        RECT 224.995 122.090 227.155 123.275 ;
        RECT 271.995 122.900 274.155 124.080 ;
        RECT 224.995 120.435 227.155 121.620 ;
        RECT 271.995 121.240 274.155 122.420 ;
        RECT 199.165 117.190 201.325 119.050 ;
        RECT 220.165 118.360 222.325 120.220 ;
        RECT 224.995 118.780 227.155 119.965 ;
        RECT 271.995 119.580 274.155 120.760 ;
        RECT 199.165 114.850 201.325 116.710 ;
        RECT 220.165 116.020 222.325 117.880 ;
        RECT 224.995 117.125 227.155 118.310 ;
        RECT 271.995 117.920 274.155 119.100 ;
        RECT 199.165 112.510 201.325 114.370 ;
        RECT 220.165 113.680 222.325 115.540 ;
        RECT 224.995 115.470 227.155 116.655 ;
        RECT 271.995 116.260 274.155 117.440 ;
        RECT 224.995 113.815 227.155 115.000 ;
        RECT 271.995 114.600 274.155 115.780 ;
        RECT 199.165 110.170 201.325 112.030 ;
        RECT 220.165 111.340 222.325 113.200 ;
        RECT 224.995 112.160 227.155 113.345 ;
        RECT 271.995 112.940 274.155 114.120 ;
        RECT 199.165 107.830 201.325 109.690 ;
        RECT 220.165 109.000 222.325 110.860 ;
        RECT 224.995 110.505 227.155 111.690 ;
        RECT 271.995 111.280 274.155 112.460 ;
        RECT 225.025 110.500 227.130 110.505 ;
        RECT 224.995 108.850 227.155 110.035 ;
        RECT 271.995 109.620 274.155 110.800 ;
        RECT 225.025 108.840 227.130 108.850 ;
        RECT 199.165 105.490 201.325 107.350 ;
        RECT 220.165 106.660 222.325 108.520 ;
        RECT 224.995 107.195 227.155 108.380 ;
        RECT 271.995 107.960 274.155 109.140 ;
        RECT 225.025 107.180 227.130 107.195 ;
        RECT 199.165 103.150 201.325 105.010 ;
        RECT 220.165 104.320 222.325 106.180 ;
        RECT 224.995 105.540 227.155 106.725 ;
        RECT 271.995 106.300 274.155 107.480 ;
        RECT 225.025 105.520 227.130 105.540 ;
        RECT 224.995 103.885 227.155 105.070 ;
        RECT 271.995 104.640 274.155 105.820 ;
        RECT 225.025 103.860 227.130 103.885 ;
        RECT 220.190 103.200 222.295 103.790 ;
        RECT 220.995 102.165 221.605 103.200 ;
        RECT 224.995 102.230 227.155 103.415 ;
        RECT 271.995 102.980 274.155 104.160 ;
        RECT 225.025 102.200 227.130 102.230 ;
        RECT 197.440 101.680 221.605 102.165 ;
        RECT 147.105 98.610 149.265 99.790 ;
        RECT 194.105 99.440 196.265 100.620 ;
        RECT 147.105 96.950 149.265 98.130 ;
        RECT 194.105 97.780 196.265 98.960 ;
        RECT 147.105 95.290 149.265 96.470 ;
        RECT 194.105 96.120 196.265 97.300 ;
        RECT 206.710 96.770 206.930 101.680 ;
        RECT 210.435 100.790 211.225 100.870 ;
        RECT 210.435 100.545 215.880 100.790 ;
        RECT 210.435 100.475 211.225 100.545 ;
        RECT 208.985 99.545 209.905 99.640 ;
        RECT 208.985 99.495 212.685 99.545 ;
        RECT 208.055 99.330 212.685 99.495 ;
        RECT 208.055 99.275 209.935 99.330 ;
        RECT 208.055 98.900 208.275 99.275 ;
        RECT 208.985 99.215 209.905 99.275 ;
        RECT 212.245 99.150 212.665 99.330 ;
        RECT 212.835 99.305 215.370 99.555 ;
        RECT 211.840 99.100 212.045 99.105 ;
        RECT 209.975 98.950 210.765 98.995 ;
        RECT 207.955 98.670 208.375 98.900 ;
        RECT 208.605 98.745 210.795 98.950 ;
        RECT 208.605 98.620 208.810 98.745 ;
        RECT 208.580 98.160 208.810 98.620 ;
        RECT 209.975 98.600 210.765 98.745 ;
        RECT 211.840 98.640 212.085 99.100 ;
        RECT 208.605 98.135 208.810 98.160 ;
        RECT 211.840 97.695 212.045 98.640 ;
        RECT 212.245 98.455 212.665 98.590 ;
        RECT 212.835 98.455 213.085 99.305 ;
        RECT 214.935 99.150 215.355 99.305 ;
        RECT 215.635 99.100 215.880 100.545 ;
        RECT 215.515 98.670 215.880 99.100 ;
        RECT 215.515 98.640 215.745 98.670 ;
        RECT 212.240 98.205 213.085 98.455 ;
        RECT 211.840 97.400 212.785 97.695 ;
        RECT 211.950 97.310 212.785 97.400 ;
        RECT 206.700 96.600 212.645 96.770 ;
        RECT 206.700 96.550 212.665 96.600 ;
        RECT 208.050 95.820 208.270 96.550 ;
        RECT 212.245 96.370 212.665 96.550 ;
        RECT 212.835 96.555 215.370 96.805 ;
        RECT 209.945 96.165 210.235 96.205 ;
        RECT 211.855 96.165 212.085 96.320 ;
        RECT 209.945 95.960 212.085 96.165 ;
        RECT 147.105 93.630 149.265 94.810 ;
        RECT 194.105 94.460 196.265 95.640 ;
        RECT 207.955 95.590 208.375 95.820 ;
        RECT 204.405 95.540 204.665 95.570 ;
        RECT 204.405 95.080 204.720 95.540 ;
        RECT 208.580 95.430 208.810 95.540 ;
        RECT 209.945 95.430 210.235 95.960 ;
        RECT 211.855 95.860 212.085 95.960 ;
        RECT 212.245 95.680 212.665 95.810 ;
        RECT 212.835 95.680 213.085 96.555 ;
        RECT 214.935 96.370 215.355 96.555 ;
        RECT 215.650 96.320 215.940 96.330 ;
        RECT 215.515 95.860 215.940 96.320 ;
        RECT 212.235 95.430 213.085 95.680 ;
        RECT 208.580 95.225 210.235 95.430 ;
        RECT 208.580 95.080 208.810 95.225 ;
        RECT 147.105 91.970 149.265 93.150 ;
        RECT 194.105 92.800 196.265 93.980 ;
        RECT 204.405 92.460 204.665 95.080 ;
        RECT 204.925 94.850 205.345 95.030 ;
        RECT 207.955 94.850 208.375 95.030 ;
        RECT 204.925 94.800 208.385 94.850 ;
        RECT 204.945 94.645 208.385 94.800 ;
        RECT 209.485 93.915 209.705 95.225 ;
        RECT 209.945 95.175 210.235 95.225 ;
        RECT 209.485 93.820 212.635 93.915 ;
        RECT 209.485 93.695 212.665 93.820 ;
        RECT 209.485 92.865 209.705 93.695 ;
        RECT 212.245 93.590 212.665 93.695 ;
        RECT 212.850 93.755 215.365 94.005 ;
        RECT 211.855 93.405 212.085 93.540 ;
        RECT 207.935 92.645 209.705 92.865 ;
        RECT 209.985 93.200 212.085 93.405 ;
        RECT 207.955 92.510 208.375 92.645 ;
        RECT 147.105 90.310 149.265 91.490 ;
        RECT 194.105 91.140 196.265 92.320 ;
        RECT 204.405 92.000 204.720 92.460 ;
        RECT 208.580 92.310 208.810 92.460 ;
        RECT 209.985 92.310 210.190 93.200 ;
        RECT 211.855 93.080 212.085 93.200 ;
        RECT 212.245 92.935 212.665 93.030 ;
        RECT 212.850 92.935 213.100 93.755 ;
        RECT 214.935 93.590 215.355 93.755 ;
        RECT 215.650 93.540 215.940 95.860 ;
        RECT 216.250 93.935 216.445 101.680 ;
        RECT 224.995 100.575 227.155 101.760 ;
        RECT 271.995 101.320 274.155 102.500 ;
        RECT 225.025 100.540 227.130 100.575 ;
        RECT 224.995 98.920 227.155 100.105 ;
        RECT 271.995 99.660 274.155 100.840 ;
        RECT 225.025 98.880 227.130 98.920 ;
        RECT 224.995 97.265 227.155 98.450 ;
        RECT 271.995 98.000 274.155 99.180 ;
        RECT 225.025 97.220 227.130 97.265 ;
        RECT 224.995 95.610 227.155 96.795 ;
        RECT 271.995 96.340 274.155 97.520 ;
        RECT 225.025 95.560 227.130 95.610 ;
        RECT 224.995 93.955 227.155 95.140 ;
        RECT 271.995 94.680 274.155 95.860 ;
        RECT 216.250 93.740 219.000 93.935 ;
        RECT 225.025 93.900 227.130 93.955 ;
        RECT 218.565 93.580 218.985 93.740 ;
        RECT 215.515 93.080 215.940 93.540 ;
        RECT 219.225 93.530 219.505 93.570 ;
        RECT 212.230 92.685 213.100 92.935 ;
        RECT 208.580 92.105 210.190 92.310 ;
        RECT 208.580 92.000 208.810 92.105 ;
        RECT 147.105 88.650 149.265 89.830 ;
        RECT 194.105 89.480 196.265 90.660 ;
        RECT 204.405 89.380 204.665 92.000 ;
        RECT 204.925 91.720 205.345 91.950 ;
        RECT 207.955 91.720 208.375 91.950 ;
        RECT 204.945 91.515 208.385 91.720 ;
        RECT 209.510 91.145 209.730 92.105 ;
        RECT 209.510 90.925 212.685 91.145 ;
        RECT 212.850 90.935 215.365 91.185 ;
        RECT 209.510 89.865 209.730 90.925 ;
        RECT 212.245 90.810 212.665 90.925 ;
        RECT 212.245 90.140 212.665 90.250 ;
        RECT 212.850 90.140 213.100 90.935 ;
        RECT 214.935 90.810 215.355 90.935 ;
        RECT 215.650 90.760 215.940 93.080 ;
        RECT 219.145 93.070 219.505 93.530 ;
        RECT 215.515 90.300 215.940 90.760 ;
        RECT 219.225 90.750 219.505 93.070 ;
        RECT 224.995 92.300 227.155 93.485 ;
        RECT 271.995 93.020 274.155 94.200 ;
        RECT 225.025 92.240 227.130 92.300 ;
        RECT 212.245 90.020 213.100 90.140 ;
        RECT 212.250 89.890 213.100 90.020 ;
        RECT 207.940 89.645 209.730 89.865 ;
        RECT 207.955 89.430 208.375 89.645 ;
        RECT 204.405 89.140 204.720 89.380 ;
        RECT 147.105 86.990 149.265 88.170 ;
        RECT 194.105 87.820 196.265 89.000 ;
        RECT 204.400 88.920 204.720 89.140 ;
        RECT 204.400 88.890 204.665 88.920 ;
        RECT 147.105 85.330 149.265 86.510 ;
        RECT 194.105 86.160 196.265 87.340 ;
        RECT 204.400 87.280 204.660 88.890 ;
        RECT 204.925 88.725 205.345 88.870 ;
        RECT 207.955 88.725 208.375 88.870 ;
        RECT 204.925 88.640 208.375 88.725 ;
        RECT 204.930 88.520 208.370 88.640 ;
        RECT 211.035 88.260 212.625 88.485 ;
        RECT 211.035 88.225 212.665 88.260 ;
        RECT 211.035 87.280 211.295 88.225 ;
        RECT 212.245 88.030 212.665 88.225 ;
        RECT 212.850 88.215 215.375 88.465 ;
        RECT 215.650 88.380 215.940 90.300 ;
        RECT 219.145 90.290 219.505 90.750 ;
        RECT 224.995 90.645 227.155 91.830 ;
        RECT 271.995 91.360 274.155 92.540 ;
        RECT 225.025 90.580 227.130 90.645 ;
        RECT 215.650 88.250 218.960 88.380 ;
        RECT 204.400 87.020 211.295 87.280 ;
        RECT 211.760 87.520 212.085 87.980 ;
        RECT 205.025 86.580 205.265 87.020 ;
        RECT 208.060 86.580 208.305 87.020 ;
        RECT 204.925 86.350 205.345 86.580 ;
        RECT 207.955 86.350 208.375 86.580 ;
        RECT 208.670 86.300 208.930 87.020 ;
        RECT 204.490 86.290 204.720 86.300 ;
        RECT 204.425 85.840 204.720 86.290 ;
        RECT 208.580 85.840 208.930 86.300 ;
        RECT 194.105 84.500 196.265 85.680 ;
        RECT 204.425 84.085 204.635 85.840 ;
        RECT 208.670 85.815 208.930 85.840 ;
        RECT 211.760 86.540 212.030 87.520 ;
        RECT 212.245 87.405 212.665 87.470 ;
        RECT 212.850 87.405 213.100 88.215 ;
        RECT 214.935 88.030 215.355 88.215 ;
        RECT 215.650 88.160 218.985 88.250 ;
        RECT 215.650 87.980 215.940 88.160 ;
        RECT 218.565 88.020 218.985 88.160 ;
        RECT 215.515 87.520 215.940 87.980 ;
        RECT 219.225 87.970 219.505 90.290 ;
        RECT 224.995 88.990 227.155 90.175 ;
        RECT 271.995 89.700 274.155 90.880 ;
        RECT 225.025 88.920 227.130 88.990 ;
        RECT 212.245 87.240 213.100 87.405 ;
        RECT 212.270 87.155 213.100 87.240 ;
        RECT 211.760 86.155 212.745 86.540 ;
        RECT 211.760 85.200 212.030 86.155 ;
        RECT 215.650 85.680 215.940 87.520 ;
        RECT 219.145 87.510 219.505 87.970 ;
        RECT 219.225 86.115 219.505 87.510 ;
        RECT 224.995 87.335 227.155 88.520 ;
        RECT 271.995 88.040 274.155 89.220 ;
        RECT 225.025 87.260 227.130 87.335 ;
        RECT 219.225 86.020 220.145 86.115 ;
        RECT 219.225 85.740 220.180 86.020 ;
        RECT 212.240 85.590 215.940 85.680 ;
        RECT 219.260 85.660 220.145 85.740 ;
        RECT 224.995 85.680 227.155 86.865 ;
        RECT 271.995 86.380 274.155 87.560 ;
        RECT 225.025 85.600 227.130 85.680 ;
        RECT 212.240 85.470 218.940 85.590 ;
        RECT 212.240 85.395 218.985 85.470 ;
        RECT 212.245 85.250 212.665 85.395 ;
        RECT 214.935 85.250 215.355 85.395 ;
        RECT 215.650 85.315 218.985 85.395 ;
        RECT 215.650 85.200 215.940 85.315 ;
        RECT 218.565 85.240 218.985 85.315 ;
        RECT 211.760 84.740 212.085 85.200 ;
        RECT 215.515 84.815 215.940 85.200 ;
        RECT 215.515 84.740 215.745 84.815 ;
        RECT 203.795 83.745 204.780 84.085 ;
        RECT 207.725 83.735 209.085 83.830 ;
        RECT 211.760 83.735 212.030 84.740 ;
        RECT 212.245 84.460 212.665 84.690 ;
        RECT 217.080 84.555 217.420 85.140 ;
        RECT 219.145 85.090 219.375 85.190 ;
        RECT 220.380 85.090 220.720 85.140 ;
        RECT 219.145 84.830 220.720 85.090 ;
        RECT 219.145 84.730 219.375 84.830 ;
        RECT 218.565 84.555 218.985 84.680 ;
        RECT 207.725 83.465 212.030 83.735 ;
        RECT 212.300 83.765 212.600 84.460 ;
        RECT 217.080 84.450 218.985 84.555 ;
        RECT 217.080 84.305 218.965 84.450 ;
        RECT 217.080 84.050 217.420 84.305 ;
        RECT 220.380 84.040 220.720 84.830 ;
        RECT 224.995 84.025 227.155 85.210 ;
        RECT 271.995 84.720 274.155 85.900 ;
        RECT 225.025 83.940 227.130 84.025 ;
        RECT 212.300 83.465 224.005 83.765 ;
        RECT 207.725 83.355 209.085 83.465 ;
        RECT 217.045 83.190 217.990 83.265 ;
        RECT 212.290 83.090 217.990 83.190 ;
        RECT 219.040 83.125 219.925 83.215 ;
        RECT 206.635 82.865 217.990 83.090 ;
        RECT 206.635 82.765 212.560 82.865 ;
        RECT 217.045 82.810 217.990 82.865 ;
        RECT 218.460 82.825 219.925 83.125 ;
        RECT 206.635 82.740 206.990 82.765 ;
        RECT 200.295 82.440 206.990 82.740 ;
        RECT 218.460 82.625 218.760 82.825 ;
        RECT 219.040 82.760 219.925 82.825 ;
        RECT 195.885 82.415 206.990 82.440 ;
        RECT 195.885 82.115 200.875 82.415 ;
        RECT 212.820 82.325 218.760 82.625 ;
        RECT 203.990 82.120 204.875 82.205 ;
        RECT 147.155 80.670 149.315 81.850 ;
        RECT 195.885 81.800 196.210 82.115 ;
        RECT 194.180 81.550 196.285 81.800 ;
        RECT 203.990 81.765 204.880 82.120 ;
        RECT 212.820 82.105 213.120 82.325 ;
        RECT 147.155 79.010 149.315 80.190 ;
        RECT 194.155 79.840 196.315 81.020 ;
        RECT 202.930 80.520 203.930 81.520 ;
        RECT 147.155 77.350 149.315 78.530 ;
        RECT 194.155 78.180 196.315 79.360 ;
        RECT 203.240 79.100 203.480 80.520 ;
        RECT 204.575 80.260 204.880 81.765 ;
        RECT 206.265 81.795 213.120 82.105 ;
        RECT 220.395 82.080 220.735 82.990 ;
        RECT 213.875 81.890 220.735 82.080 ;
        RECT 206.265 81.520 206.575 81.795 ;
        RECT 213.875 81.780 220.730 81.890 ;
        RECT 205.620 80.520 206.620 81.520 ;
        RECT 213.875 81.490 214.175 81.780 ;
        RECT 203.990 79.955 204.880 80.260 ;
        RECT 201.090 78.880 201.320 79.010 ;
        RECT 202.060 78.880 202.290 79.010 ;
        RECT 203.200 78.880 203.530 79.100 ;
        RECT 201.090 78.680 203.530 78.880 ;
        RECT 201.090 78.550 201.320 78.680 ;
        RECT 202.060 78.550 202.290 78.680 ;
        RECT 203.200 78.510 203.530 78.680 ;
        RECT 201.480 78.310 201.900 78.500 ;
        RECT 203.990 78.310 204.295 79.955 ;
        RECT 206.250 79.790 206.580 80.520 ;
        RECT 207.360 80.490 208.360 81.490 ;
        RECT 213.220 80.490 214.220 81.490 ;
        RECT 214.960 80.520 215.960 81.520 ;
        RECT 217.650 80.520 218.650 81.520 ;
        RECT 207.400 79.790 207.730 80.490 ;
        RECT 213.850 79.790 214.180 80.490 ;
        RECT 215.000 79.790 215.330 80.520 ;
        RECT 204.980 79.300 208.740 79.590 ;
        RECT 212.840 79.300 216.600 79.590 ;
        RECT 204.975 79.260 208.745 79.300 ;
        RECT 204.490 78.860 204.820 79.090 ;
        RECT 204.975 79.070 205.395 79.260 ;
        RECT 208.325 79.070 208.745 79.260 ;
        RECT 212.835 79.260 216.605 79.300 ;
        RECT 212.835 79.070 213.255 79.260 ;
        RECT 216.185 79.070 216.605 79.260 ;
        RECT 218.100 79.100 218.340 80.520 ;
        RECT 205.600 78.860 205.830 79.020 ;
        RECT 207.890 78.930 208.120 79.020 ;
        RECT 208.950 78.930 209.180 79.020 ;
        RECT 204.490 78.650 205.910 78.860 ;
        RECT 207.390 78.670 209.180 78.930 ;
        RECT 204.490 78.500 204.820 78.650 ;
        RECT 205.600 78.560 205.830 78.650 ;
        RECT 204.975 78.310 205.395 78.510 ;
        RECT 207.390 78.380 207.650 78.670 ;
        RECT 207.890 78.560 208.120 78.670 ;
        RECT 208.950 78.560 209.180 78.670 ;
        RECT 212.400 78.930 212.630 79.020 ;
        RECT 213.460 78.930 213.690 79.020 ;
        RECT 212.400 78.670 214.190 78.930 ;
        RECT 215.750 78.860 215.980 79.020 ;
        RECT 216.760 78.860 217.090 79.090 ;
        RECT 212.400 78.560 212.630 78.670 ;
        RECT 213.460 78.560 213.690 78.670 ;
        RECT 213.930 78.380 214.190 78.670 ;
        RECT 215.670 78.650 217.090 78.860 ;
        RECT 215.750 78.560 215.980 78.650 ;
        RECT 205.580 78.310 205.910 78.380 ;
        RECT 207.360 78.310 207.690 78.380 ;
        RECT 201.440 78.050 207.690 78.310 ;
        RECT 205.580 77.790 205.910 78.050 ;
        RECT 207.360 77.790 207.690 78.050 ;
        RECT 213.890 78.310 214.220 78.380 ;
        RECT 215.670 78.310 216.000 78.380 ;
        RECT 216.185 78.310 216.605 78.510 ;
        RECT 216.760 78.500 217.090 78.650 ;
        RECT 218.050 78.880 218.380 79.100 ;
        RECT 219.290 78.880 219.520 79.010 ;
        RECT 220.260 78.880 220.490 79.010 ;
        RECT 218.050 78.680 220.490 78.880 ;
        RECT 218.050 78.510 218.380 78.680 ;
        RECT 219.290 78.550 219.520 78.680 ;
        RECT 220.260 78.550 220.490 78.680 ;
        RECT 219.680 78.310 220.100 78.500 ;
        RECT 213.890 78.050 220.140 78.310 ;
        RECT 213.890 77.790 214.220 78.050 ;
        RECT 215.670 77.790 216.000 78.050 ;
        RECT 147.155 75.690 149.315 76.870 ;
        RECT 194.155 76.520 196.315 77.700 ;
        RECT 204.490 76.460 204.820 76.740 ;
        RECT 206.240 76.460 206.570 76.730 ;
        RECT 215.010 76.460 215.340 76.730 ;
        RECT 216.760 76.460 217.090 76.740 ;
        RECT 201.460 76.200 207.660 76.460 ;
        RECT 147.155 74.030 149.315 75.210 ;
        RECT 194.155 74.860 196.315 76.040 ;
        RECT 201.470 76.030 201.890 76.200 ;
        RECT 204.490 76.150 204.820 76.200 ;
        RECT 204.985 76.020 205.405 76.200 ;
        RECT 206.240 76.140 206.570 76.200 ;
        RECT 204.550 75.860 204.780 75.970 ;
        RECT 205.590 75.860 205.920 76.040 ;
        RECT 204.550 75.650 205.920 75.860 ;
        RECT 204.550 75.510 204.780 75.650 ;
        RECT 204.985 75.250 205.405 75.460 ;
        RECT 205.590 75.450 205.920 75.650 ;
        RECT 207.400 75.840 207.660 76.200 ;
        RECT 213.920 76.200 220.120 76.460 ;
        RECT 207.890 75.840 208.120 75.940 ;
        RECT 208.950 75.840 209.180 75.940 ;
        RECT 207.400 75.580 209.180 75.840 ;
        RECT 207.890 75.480 208.120 75.580 ;
        RECT 208.950 75.480 209.180 75.580 ;
        RECT 212.400 75.840 212.630 75.940 ;
        RECT 213.460 75.840 213.690 75.940 ;
        RECT 213.920 75.840 214.180 76.200 ;
        RECT 215.010 76.140 215.340 76.200 ;
        RECT 212.400 75.580 214.180 75.840 ;
        RECT 215.660 75.860 215.990 76.040 ;
        RECT 216.175 76.020 216.595 76.200 ;
        RECT 216.760 76.150 217.090 76.200 ;
        RECT 219.690 76.030 220.110 76.200 ;
        RECT 216.800 75.860 217.030 75.970 ;
        RECT 215.660 75.650 217.030 75.860 ;
        RECT 212.400 75.480 212.630 75.580 ;
        RECT 213.460 75.480 213.690 75.580 ;
        RECT 215.660 75.450 215.990 75.650 ;
        RECT 216.800 75.510 217.030 75.650 ;
        RECT 208.325 75.250 208.745 75.430 ;
        RECT 204.980 75.200 208.745 75.250 ;
        RECT 212.835 75.250 213.255 75.430 ;
        RECT 216.175 75.250 216.595 75.460 ;
        RECT 212.835 75.200 216.600 75.250 ;
        RECT 204.980 74.920 208.740 75.200 ;
        RECT 212.840 74.920 216.600 75.200 ;
        RECT 147.155 72.370 149.315 73.550 ;
        RECT 194.155 73.200 196.315 74.380 ;
        RECT 147.155 70.710 149.315 71.890 ;
        RECT 194.155 71.540 196.315 72.720 ;
        RECT 147.155 69.050 149.315 70.230 ;
        RECT 194.155 69.880 196.315 71.060 ;
        RECT 215.820 70.920 217.925 70.960 ;
        RECT 215.820 70.430 221.805 70.920 ;
        RECT 215.820 70.370 217.925 70.430 ;
        RECT 147.155 67.390 149.315 68.570 ;
        RECT 194.155 68.220 196.315 69.400 ;
        RECT 203.200 67.970 203.530 68.460 ;
        RECT 209.615 68.110 209.875 68.660 ;
        RECT 203.170 67.810 207.020 67.970 ;
        RECT 202.800 67.760 207.020 67.810 ;
        RECT 194.155 66.560 196.315 67.740 ;
        RECT 202.800 67.580 203.800 67.760 ;
        RECT 205.990 67.580 206.990 67.760 ;
        RECT 209.620 67.195 209.820 68.110 ;
        RECT 218.050 67.970 218.380 68.460 ;
        RECT 214.560 67.810 218.410 67.970 ;
        RECT 214.560 67.760 218.780 67.810 ;
        RECT 214.590 67.580 215.590 67.760 ;
        RECT 217.780 67.580 218.780 67.760 ;
        RECT 209.620 67.160 209.855 67.195 ;
        RECT 208.720 66.950 209.855 67.160 ;
        RECT 206.880 65.075 207.110 65.130 ;
        RECT 208.720 65.075 208.920 66.950 ;
        RECT 209.625 66.905 209.855 66.950 ;
        RECT 210.015 66.715 210.515 66.945 ;
        RECT 210.110 65.320 210.335 66.715 ;
        RECT 211.895 66.405 212.170 66.775 ;
        RECT 210.015 65.090 210.515 65.320 ;
        RECT 211.945 65.130 212.115 66.405 ;
        RECT 221.315 65.765 221.805 70.430 ;
        RECT 223.705 66.810 224.005 83.465 ;
        RECT 224.995 82.370 227.155 83.555 ;
        RECT 271.995 83.060 274.155 84.240 ;
        RECT 225.025 82.280 227.130 82.370 ;
        RECT 224.995 80.715 227.155 81.900 ;
        RECT 271.995 81.400 274.155 82.580 ;
        RECT 225.025 80.620 227.130 80.715 ;
        RECT 224.995 79.060 227.155 80.245 ;
        RECT 271.995 79.740 274.155 80.920 ;
        RECT 225.025 78.960 227.130 79.060 ;
        RECT 224.995 77.405 227.155 78.590 ;
        RECT 271.995 78.080 274.155 79.260 ;
        RECT 225.025 77.300 227.130 77.405 ;
        RECT 224.995 75.750 227.155 76.935 ;
        RECT 271.995 76.420 274.155 77.600 ;
        RECT 225.025 75.640 227.130 75.750 ;
        RECT 224.995 74.095 227.155 75.280 ;
        RECT 271.995 74.760 274.155 75.940 ;
        RECT 225.025 73.980 227.130 74.095 ;
        RECT 224.995 72.440 227.155 73.625 ;
        RECT 271.995 73.100 274.155 74.280 ;
        RECT 225.025 72.320 227.130 72.440 ;
        RECT 224.995 70.785 227.155 71.970 ;
        RECT 271.995 71.440 274.155 72.620 ;
        RECT 225.025 70.660 227.130 70.785 ;
        RECT 224.995 69.130 227.155 70.315 ;
        RECT 271.995 69.780 274.155 70.960 ;
        RECT 225.025 69.000 227.130 69.130 ;
        RECT 224.995 67.475 227.155 68.660 ;
        RECT 271.995 68.120 274.155 69.300 ;
        RECT 225.025 67.340 227.130 67.475 ;
        RECT 223.705 66.460 227.155 66.810 ;
        RECT 271.995 66.460 274.155 67.640 ;
        RECT 212.925 65.275 221.805 65.765 ;
        RECT 205.675 64.690 206.675 64.880 ;
        RECT 206.880 64.875 208.920 65.075 ;
        RECT 206.880 64.840 207.110 64.875 ;
        RECT 210.015 64.690 210.515 64.880 ;
        RECT 211.915 64.840 212.145 65.130 ;
        RECT 212.305 64.690 212.725 64.880 ;
        RECT 212.925 64.690 213.415 65.275 ;
        RECT 205.660 64.195 213.415 64.690 ;
      LAYER via ;
        RECT 210.540 100.545 210.800 100.805 ;
        RECT 210.860 100.545 211.120 100.805 ;
        RECT 208.995 99.300 209.255 99.560 ;
        RECT 209.315 99.300 209.575 99.560 ;
        RECT 209.635 99.300 209.895 99.560 ;
        RECT 210.080 98.670 210.340 98.930 ;
        RECT 210.400 98.670 210.660 98.930 ;
        RECT 212.080 97.375 212.340 97.635 ;
        RECT 212.400 97.375 212.660 97.635 ;
        RECT 209.960 95.880 210.220 96.140 ;
        RECT 209.960 95.560 210.220 95.820 ;
        RECT 209.960 95.240 210.220 95.500 ;
        RECT 212.040 86.220 212.300 86.480 ;
        RECT 212.360 86.220 212.620 86.480 ;
        RECT 219.415 85.760 219.675 86.020 ;
        RECT 219.735 85.760 219.995 86.020 ;
        RECT 217.120 84.790 217.380 85.050 ;
        RECT 204.000 83.785 204.260 84.045 ;
        RECT 204.320 83.785 204.580 84.045 ;
        RECT 220.420 84.780 220.680 85.040 ;
        RECT 217.120 84.470 217.380 84.730 ;
        RECT 207.795 83.465 208.055 83.725 ;
        RECT 208.115 83.465 208.375 83.725 ;
        RECT 208.435 83.465 208.695 83.725 ;
        RECT 208.755 83.465 209.015 83.725 ;
        RECT 220.420 84.460 220.680 84.720 ;
        RECT 217.120 84.150 217.380 84.410 ;
        RECT 220.420 84.140 220.680 84.400 ;
        RECT 217.260 82.910 217.520 83.170 ;
        RECT 217.580 82.910 217.840 83.170 ;
        RECT 219.195 82.860 219.455 83.120 ;
        RECT 219.515 82.860 219.775 83.120 ;
        RECT 220.435 82.630 220.695 82.890 ;
        RECT 204.145 81.855 204.405 82.115 ;
        RECT 204.465 81.855 204.725 82.115 ;
        RECT 220.435 82.310 220.695 82.570 ;
        RECT 220.435 81.990 220.695 82.250 ;
        RECT 206.285 79.955 206.545 80.215 ;
        RECT 203.235 78.675 203.495 78.935 ;
        RECT 207.435 79.955 207.695 80.215 ;
        RECT 213.885 79.955 214.145 80.215 ;
        RECT 215.035 79.955 215.295 80.215 ;
        RECT 204.525 78.665 204.785 78.925 ;
        RECT 216.795 78.665 217.055 78.925 ;
        RECT 205.615 77.955 205.875 78.215 ;
        RECT 207.395 77.955 207.655 78.215 ;
        RECT 218.085 78.675 218.345 78.935 ;
        RECT 213.925 77.955 214.185 78.215 ;
        RECT 215.705 77.955 215.965 78.215 ;
        RECT 204.525 76.315 204.785 76.575 ;
        RECT 206.275 76.305 206.535 76.565 ;
        RECT 205.625 75.615 205.885 75.875 ;
        RECT 215.045 76.305 215.305 76.565 ;
        RECT 216.795 76.315 217.055 76.575 ;
        RECT 215.695 75.615 215.955 75.875 ;
        RECT 203.235 68.035 203.495 68.295 ;
        RECT 209.615 68.255 209.875 68.515 ;
        RECT 218.085 68.035 218.345 68.295 ;
        RECT 211.905 66.460 212.165 66.720 ;
      LAYER met2 ;
        RECT 210.385 100.525 211.275 100.820 ;
        RECT 208.935 99.265 209.955 99.590 ;
        RECT 209.310 85.080 209.570 99.265 ;
        RECT 210.455 98.945 210.680 100.525 ;
        RECT 209.925 98.650 210.815 98.945 ;
        RECT 209.985 96.155 210.210 98.650 ;
        RECT 211.900 97.360 212.835 97.645 ;
        RECT 209.895 95.225 210.285 96.155 ;
        RECT 211.995 86.490 212.300 97.360 ;
        RECT 211.860 86.205 212.795 86.490 ;
        RECT 219.210 85.710 220.195 86.065 ;
        RECT 209.310 84.820 210.280 85.080 ;
        RECT 203.845 83.780 204.780 84.135 ;
        RECT 203.845 83.695 209.135 83.780 ;
        RECT 204.330 83.410 209.135 83.695 ;
        RECT 204.330 82.155 204.765 83.410 ;
        RECT 207.695 83.405 209.135 83.410 ;
        RECT 203.940 81.815 204.925 82.155 ;
        RECT 206.200 79.840 206.630 80.330 ;
        RECT 207.350 79.840 207.780 80.330 ;
        RECT 203.150 78.560 203.580 79.050 ;
        RECT 203.230 69.000 203.500 78.560 ;
        RECT 204.440 78.550 204.870 79.040 ;
        RECT 204.540 76.690 204.810 78.550 ;
        RECT 205.610 78.330 205.880 78.400 ;
        RECT 205.530 77.840 205.960 78.330 ;
        RECT 204.440 76.200 204.870 76.690 ;
        RECT 204.540 76.100 204.810 76.200 ;
        RECT 205.610 75.990 205.880 77.840 ;
        RECT 206.260 76.680 206.540 79.840 ;
        RECT 207.420 78.330 207.690 79.840 ;
        RECT 207.310 77.840 207.740 78.330 ;
        RECT 206.190 76.190 206.620 76.680 ;
        RECT 205.540 75.500 205.970 75.990 ;
        RECT 210.020 72.155 210.280 84.820 ;
        RECT 217.030 84.100 217.470 85.100 ;
        RECT 217.055 83.215 217.420 84.100 ;
        RECT 217.045 82.860 218.045 83.215 ;
        RECT 219.395 83.165 219.705 85.710 ;
        RECT 220.330 84.090 220.770 85.090 ;
        RECT 218.990 82.810 219.975 83.165 ;
        RECT 220.415 82.940 220.705 84.090 ;
        RECT 220.345 81.940 220.785 82.940 ;
        RECT 213.800 79.840 214.230 80.330 ;
        RECT 214.950 79.840 215.380 80.330 ;
        RECT 213.890 78.330 214.160 79.840 ;
        RECT 213.840 77.840 214.270 78.330 ;
        RECT 215.040 76.680 215.320 79.840 ;
        RECT 216.710 78.550 217.140 79.040 ;
        RECT 218.000 78.560 218.430 79.050 ;
        RECT 215.700 78.330 215.970 78.400 ;
        RECT 215.620 77.840 216.050 78.330 ;
        RECT 214.960 76.190 215.390 76.680 ;
        RECT 215.700 75.990 215.970 77.840 ;
        RECT 216.770 76.690 217.040 78.550 ;
        RECT 216.710 76.200 217.140 76.690 ;
        RECT 216.770 76.100 217.040 76.200 ;
        RECT 215.610 75.500 216.040 75.990 ;
        RECT 209.620 71.895 210.280 72.155 ;
        RECT 203.230 68.410 203.545 69.000 ;
        RECT 209.620 68.610 209.880 71.895 ;
        RECT 203.150 67.920 203.580 68.410 ;
        RECT 209.565 68.160 209.920 68.610 ;
        RECT 218.080 68.410 218.350 78.560 ;
        RECT 218.000 67.920 218.430 68.410 ;
        RECT 203.275 66.725 203.545 67.920 ;
        RECT 203.275 66.455 212.235 66.725 ;
  END
END sky130_ef_ip__xtal_osc_32k_DI
END LIBRARY

