magic
tech sky130A
magscale 1 2
timestamp 1527799877
<< checkpaint >>
rect 11751 -1916 116199 44965
<< via1 >>
rect 40723 26665 40839 26781
rect 51601 12831 51717 12947
<< metal2 >>
rect 13011 28464 13139 43705
rect 114811 33393 114939 43705
rect 55850 33173 114939 33393
rect 13011 28216 40880 28464
rect 40680 26781 40880 28216
rect 40680 26665 40723 26781
rect 40839 26665 40880 26781
rect 40680 26620 40880 26665
tri 40880 26658 40881 28464 nw
rect 55850 26620 56050 33173
rect 51562 12947 51762 12986
rect 51562 12831 51601 12947
rect 51717 12831 51762 12947
rect 51562 0 51762 12831
rect 52402 0 52602 12863
rect 54885 0 55085 12863
rect 51562 -656 51618 0
rect 52402 -656 52458 0
rect 54885 -656 54941 0
<< via2 >>
rect 42915 26513 43211 26800
rect 43581 26513 43877 26800
rect 44240 26509 44536 26796
rect 44903 26509 45199 26796
rect 47044 26513 47340 26800
rect 47710 26513 48006 26800
rect 48369 26509 48665 26796
rect 49032 26509 49328 26796
rect 58352 26513 58648 26800
rect 59018 26513 59314 26800
rect 59677 26509 59973 26796
rect 60340 26509 60636 26796
rect 62481 26513 62777 26800
rect 63147 26513 63443 26800
rect 63806 26509 64102 26796
rect 64469 26509 64765 26796
rect 42915 12821 43211 13108
rect 43581 12821 43877 13108
rect 44240 12817 44536 13104
rect 44903 12817 45199 13104
rect 47044 12821 47340 13108
rect 47710 12821 48006 13108
rect 48369 12817 48665 13104
rect 49032 12817 49328 13104
rect 51965 12860 52101 13620
rect 54440 12860 54576 13564
rect 58352 12821 58648 13108
rect 59018 12821 59314 13108
rect 59677 12817 59973 13104
rect 60340 12817 60636 13104
rect 62481 12821 62777 13108
rect 63147 12821 63443 13108
rect 63806 12817 64102 13104
rect 64469 12817 64765 13104
<< metal3 >>
rect 41866 26804 45866 26820
rect 41866 26509 42911 26804
rect 43215 26509 43577 26804
rect 43881 26800 45866 26804
rect 43881 26509 44236 26800
rect 41866 26505 44236 26509
rect 44540 26505 44899 26800
rect 45203 26505 45866 26800
rect 41866 26478 45866 26505
rect 46151 26804 50151 26820
rect 46151 26509 47040 26804
rect 47344 26509 47706 26804
rect 48010 26800 50151 26804
rect 48010 26509 48365 26800
rect 46151 26505 48365 26509
rect 48669 26505 49028 26800
rect 49332 26505 50151 26800
rect 46151 26478 50151 26505
rect 57303 26804 61303 26820
rect 57303 26509 58348 26804
rect 58652 26509 59014 26804
rect 59318 26800 61303 26804
rect 59318 26509 59673 26800
rect 57303 26505 59673 26509
rect 59977 26505 60336 26800
rect 60640 26505 61303 26800
rect 57303 26478 61303 26505
rect 61588 26804 65588 26820
rect 61588 26509 62477 26804
rect 62781 26509 63143 26804
rect 63447 26800 65588 26804
rect 63447 26509 63802 26800
rect 61588 26505 63802 26509
rect 64106 26505 64465 26800
rect 64769 26505 65588 26800
rect 61588 26478 65588 26505
rect 51925 13624 52125 13718
rect 41866 13112 45866 13128
rect 41866 12817 42911 13112
rect 43215 12817 43577 13112
rect 43881 13108 45866 13112
rect 43881 12817 44236 13108
rect 41866 12813 44236 12817
rect 44540 12813 44899 13108
rect 45203 12813 45866 13108
rect 41866 12786 45866 12813
rect 46151 13112 50151 13128
rect 46151 12817 47040 13112
rect 47344 12817 47706 13112
rect 48010 13108 50151 13112
rect 48010 12817 48365 13108
rect 46151 12813 48365 12817
rect 48669 12813 49028 13108
rect 49332 12813 50151 13108
rect 46151 12786 50151 12813
rect 51925 12856 51961 13624
rect 52105 12856 52125 13624
rect 51925 12786 52125 12856
rect 54400 13568 54600 13575
rect 54400 12856 54436 13568
rect 54580 12856 54600 13568
rect 54400 12786 54600 12856
rect 57303 13112 61303 13128
rect 57303 12817 58348 13112
rect 58652 12817 59014 13112
rect 59318 13108 61303 13112
rect 59318 12817 59673 13108
rect 57303 12813 59673 12817
rect 59977 12813 60336 13108
rect 60640 12813 61303 13108
rect 57303 12786 61303 12813
rect 61588 13112 65588 13128
rect 61588 12817 62477 13112
rect 62781 12817 63143 13112
rect 63447 13108 65588 13112
rect 63447 12817 63802 13108
rect 61588 12813 63802 12817
rect 64106 12813 64465 13108
rect 64769 12813 65588 13108
rect 61588 12786 65588 12813
<< via3 >>
rect 42911 26800 43215 26804
rect 42911 26513 42915 26800
rect 42915 26513 43211 26800
rect 43211 26513 43215 26800
rect 42911 26509 43215 26513
rect 43577 26800 43881 26804
rect 43577 26513 43581 26800
rect 43581 26513 43877 26800
rect 43877 26513 43881 26800
rect 43577 26509 43881 26513
rect 44236 26796 44540 26800
rect 44236 26509 44240 26796
rect 44240 26509 44536 26796
rect 44536 26509 44540 26796
rect 44236 26505 44540 26509
rect 44899 26796 45203 26800
rect 44899 26509 44903 26796
rect 44903 26509 45199 26796
rect 45199 26509 45203 26796
rect 44899 26505 45203 26509
rect 47040 26800 47344 26804
rect 47040 26513 47044 26800
rect 47044 26513 47340 26800
rect 47340 26513 47344 26800
rect 47040 26509 47344 26513
rect 47706 26800 48010 26804
rect 47706 26513 47710 26800
rect 47710 26513 48006 26800
rect 48006 26513 48010 26800
rect 47706 26509 48010 26513
rect 48365 26796 48669 26800
rect 48365 26509 48369 26796
rect 48369 26509 48665 26796
rect 48665 26509 48669 26796
rect 48365 26505 48669 26509
rect 49028 26796 49332 26800
rect 49028 26509 49032 26796
rect 49032 26509 49328 26796
rect 49328 26509 49332 26796
rect 49028 26505 49332 26509
rect 58348 26800 58652 26804
rect 58348 26513 58352 26800
rect 58352 26513 58648 26800
rect 58648 26513 58652 26800
rect 58348 26509 58652 26513
rect 59014 26800 59318 26804
rect 59014 26513 59018 26800
rect 59018 26513 59314 26800
rect 59314 26513 59318 26800
rect 59014 26509 59318 26513
rect 59673 26796 59977 26800
rect 59673 26509 59677 26796
rect 59677 26509 59973 26796
rect 59973 26509 59977 26796
rect 59673 26505 59977 26509
rect 60336 26796 60640 26800
rect 60336 26509 60340 26796
rect 60340 26509 60636 26796
rect 60636 26509 60640 26796
rect 60336 26505 60640 26509
rect 62477 26800 62781 26804
rect 62477 26513 62481 26800
rect 62481 26513 62777 26800
rect 62777 26513 62781 26800
rect 62477 26509 62781 26513
rect 63143 26800 63447 26804
rect 63143 26513 63147 26800
rect 63147 26513 63443 26800
rect 63443 26513 63447 26800
rect 63143 26509 63447 26513
rect 63802 26796 64106 26800
rect 63802 26509 63806 26796
rect 63806 26509 64102 26796
rect 64102 26509 64106 26796
rect 63802 26505 64106 26509
rect 64465 26796 64769 26800
rect 64465 26509 64469 26796
rect 64469 26509 64765 26796
rect 64765 26509 64769 26796
rect 64465 26505 64769 26509
rect 42911 13108 43215 13112
rect 42911 12821 42915 13108
rect 42915 12821 43211 13108
rect 43211 12821 43215 13108
rect 42911 12817 43215 12821
rect 43577 13108 43881 13112
rect 43577 12821 43581 13108
rect 43581 12821 43877 13108
rect 43877 12821 43881 13108
rect 43577 12817 43881 12821
rect 44236 13104 44540 13108
rect 44236 12817 44240 13104
rect 44240 12817 44536 13104
rect 44536 12817 44540 13104
rect 44236 12813 44540 12817
rect 44899 13104 45203 13108
rect 44899 12817 44903 13104
rect 44903 12817 45199 13104
rect 45199 12817 45203 13104
rect 44899 12813 45203 12817
rect 47040 13108 47344 13112
rect 47040 12821 47044 13108
rect 47044 12821 47340 13108
rect 47340 12821 47344 13108
rect 47040 12817 47344 12821
rect 47706 13108 48010 13112
rect 47706 12821 47710 13108
rect 47710 12821 48006 13108
rect 48006 12821 48010 13108
rect 47706 12817 48010 12821
rect 48365 13104 48669 13108
rect 48365 12817 48369 13104
rect 48369 12817 48665 13104
rect 48665 12817 48669 13104
rect 48365 12813 48669 12817
rect 49028 13104 49332 13108
rect 49028 12817 49032 13104
rect 49032 12817 49328 13104
rect 49328 12817 49332 13104
rect 49028 12813 49332 12817
rect 51961 13620 52105 13624
rect 51961 12860 51965 13620
rect 51965 12860 52101 13620
rect 52101 12860 52105 13620
rect 51961 12856 52105 12860
rect 54436 13564 54580 13568
rect 54436 12860 54440 13564
rect 54440 12860 54576 13564
rect 54576 12860 54580 13564
rect 54436 12856 54580 12860
rect 58348 13108 58652 13112
rect 58348 12821 58352 13108
rect 58352 12821 58648 13108
rect 58648 12821 58652 13108
rect 58348 12817 58652 12821
rect 59014 13108 59318 13112
rect 59014 12821 59018 13108
rect 59018 12821 59314 13108
rect 59314 12821 59318 13108
rect 59014 12817 59318 12821
rect 59673 13104 59977 13108
rect 59673 12817 59677 13104
rect 59677 12817 59973 13104
rect 59973 12817 59977 13104
rect 59673 12813 59977 12817
rect 60336 13104 60640 13108
rect 60336 12817 60340 13104
rect 60340 12817 60636 13104
rect 60636 12817 60640 13104
rect 60336 12813 60640 12817
rect 62477 13108 62781 13112
rect 62477 12821 62481 13108
rect 62481 12821 62777 13108
rect 62777 12821 62781 13108
rect 62477 12817 62781 12821
rect 63143 13108 63447 13112
rect 63143 12821 63147 13108
rect 63147 12821 63443 13108
rect 63443 12821 63447 13108
rect 63143 12817 63447 12821
rect 63802 13104 64106 13108
rect 63802 12817 63806 13104
rect 63806 12817 64102 13104
rect 64102 12817 64106 13104
rect 63802 12813 64106 12817
rect 64465 13104 64769 13108
rect 64465 12817 64469 13104
rect 64469 12817 64765 13104
rect 64765 12817 64769 13104
rect 64465 12813 64769 12817
<< metal4 >>
rect 42909 26804 43229 42360
rect 42909 26509 42911 26804
rect 43215 26509 43229 26804
rect 42909 13112 43229 26509
rect 42909 12817 42911 13112
rect 43215 12817 43229 13112
rect 42909 660 43229 12817
rect 43569 26804 43889 42360
rect 43569 26509 43577 26804
rect 43881 26509 43889 26804
rect 43569 13112 43889 26509
rect 43569 12817 43577 13112
rect 43881 12817 43889 13112
rect 43569 660 43889 12817
rect 44229 26800 44549 42360
rect 44229 26505 44236 26800
rect 44540 26505 44549 26800
rect 44229 13108 44549 26505
rect 44229 12813 44236 13108
rect 44540 12813 44549 13108
rect 44229 660 44549 12813
rect 44889 26800 45209 42360
rect 44889 26505 44899 26800
rect 45203 26505 45209 26800
rect 44889 13108 45209 26505
rect 44889 12813 44899 13108
rect 45203 12813 45209 13108
rect 44889 660 45209 12813
rect 47033 26804 47353 42360
rect 47033 26509 47040 26804
rect 47344 26509 47353 26804
rect 47033 13112 47353 26509
rect 47033 12817 47040 13112
rect 47344 12817 47353 13112
rect 47033 660 47353 12817
rect 47693 26804 48013 42360
rect 47693 26509 47706 26804
rect 48010 26509 48013 26804
rect 47693 13112 48013 26509
rect 47693 12817 47706 13112
rect 48010 12817 48013 13112
rect 47693 660 48013 12817
rect 48353 26800 48673 42360
rect 48353 26505 48365 26800
rect 48669 26505 48673 26800
rect 48353 13108 48673 26505
rect 48353 12813 48365 13108
rect 48669 12813 48673 13108
rect 48353 660 48673 12813
rect 49013 26800 49333 42360
rect 49013 26505 49028 26800
rect 49332 26505 49333 26800
rect 49013 13108 49333 26505
rect 49013 12813 49028 13108
rect 49332 12813 49333 13108
rect 49013 660 49333 12813
rect 51867 13624 52187 42360
rect 51867 12856 51961 13624
rect 52105 12856 52187 13624
rect 51867 660 52187 12856
rect 54334 13568 54654 42360
rect 54334 12856 54436 13568
rect 54580 12856 54654 13568
rect 54334 660 54654 12856
rect 58346 26804 58666 42360
rect 58346 26509 58348 26804
rect 58652 26509 58666 26804
rect 58346 13112 58666 26509
rect 58346 12817 58348 13112
rect 58652 12817 58666 13112
rect 58346 660 58666 12817
rect 59006 26804 59326 42360
rect 59006 26509 59014 26804
rect 59318 26509 59326 26804
rect 59006 13112 59326 26509
rect 59006 12817 59014 13112
rect 59318 12817 59326 13112
rect 59006 660 59326 12817
rect 59666 26800 59986 42360
rect 59666 26505 59673 26800
rect 59977 26505 59986 26800
rect 59666 13108 59986 26505
rect 59666 12813 59673 13108
rect 59977 12813 59986 13108
rect 59666 660 59986 12813
rect 60326 26800 60646 42360
rect 60326 26505 60336 26800
rect 60640 26505 60646 26800
rect 60326 13108 60646 26505
rect 60326 12813 60336 13108
rect 60640 12813 60646 13108
rect 60326 660 60646 12813
rect 62470 26804 62790 42360
rect 62470 26509 62477 26804
rect 62781 26509 62790 26804
rect 62470 13112 62790 26509
rect 62470 12817 62477 13112
rect 62781 12817 62790 13112
rect 62470 660 62790 12817
rect 63130 26804 63450 42360
rect 63130 26509 63143 26804
rect 63447 26509 63450 26804
rect 63130 13112 63450 26509
rect 63130 12817 63143 13112
rect 63447 12817 63450 13112
rect 63130 660 63450 12817
rect 63790 26800 64110 42360
rect 63790 26505 63802 26800
rect 64106 26505 64110 26800
rect 63790 13108 64110 26505
rect 63790 12813 63802 13108
rect 64106 12813 64110 13108
rect 63790 660 64110 12813
rect 64450 26800 64770 42360
rect 64450 26505 64465 26800
rect 64769 26505 64770 26800
rect 64450 13108 64770 26505
rect 64450 12813 64465 13108
rect 64769 12813 64770 13108
rect 64450 660 64770 12813
use sky130_ef_ip__xtal_osc_32k  mprj
timestamp 1527799877
transform 0 -1 67059 -1 0 26820
box 0 0 14034 26558
<< labels >>
flabel metal2 s 13011 42249 13139 43705 0 FreeSans 280 90 0 0 in
port 4 nsew
flabel metal2 s 114811 42249 114939 43705 0 FreeSans 280 90 0 0 out
port 3 nsew
flabel metal2 s 54885 -656 54941 144 0 FreeSans 280 90 0 0 boost
port 1 nsew
flabel metal2 s 52402 -656 52458 144 0 FreeSans 280 90 0 0 ena
port 2 nsew
flabel metal2 s 51562 -656 51618 144 0 FreeSans 280 90 0 0 dout
port 5 nsew
flabel metal4 s 44889 660 45209 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 43569 660 43889 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 42909 660 43229 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 44229 660 44549 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 49013 660 49333 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 47693 660 48013 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 47033 660 47353 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 48353 660 48673 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 60326 660 60646 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 59006 660 59326 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 59666 660 59986 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 63130 660 63450 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 62470 660 62790 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 63790 660 64110 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 51867 660 52187 42360 0 FreeSans 2400 90 0 0 vssd1
port 8 nsew
flabel metal4 s 54334 660 54654 42360 0 FreeSans 2400 90 0 0 vccd1
port 9 nsew
flabel metal4 s 64450 660 64770 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 58346 660 58666 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
<< properties >>
string FIXED_BBOX 11646 0 116706 42360
<< end >>
