VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_32k_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_32k_DI ;
  ORIGIN 0.000 0.000 ;
  SIZE 525.300 BY 211.800 ;
  PIN boost
    ANTENNAGATEAREA 0.510000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 216.195 -3.280 216.475 64.930 ;
    END
  END boost
  PIN ena
    ANTENNAGATEAREA 0.585000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 203.780 -3.280 204.060 64.930 ;
    END
  END ena
  PIN out
    PORT
      LAYER met2 ;
        RECT 515.825 165.865 516.465 218.525 ;
    END
  END out
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER met2 ;
        RECT 6.825 142.320 7.465 218.525 ;
    END
  END in
  PIN dout
    PORT
      LAYER met2 ;
        RECT 199.580 -3.280 199.860 64.155 ;
    END
  END dout
  PIN vdda1
    ANTENNADIFFAREA 200.228592 ;
    PORT
      LAYER met4 ;
        RECT 186.835 3.300 188.435 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.235 3.300 181.835 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 176.935 3.300 178.535 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.535 3.300 185.135 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 257.420 3.300 259.020 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.120 3.300 255.720 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.720 3.300 262.320 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.020 3.300 265.620 211.800 ;
    END
  END vdda1
  PIN vssa1
    ANTENNADIFFAREA 167.107590 ;
    PORT
      LAYER met4 ;
        RECT 166.215 3.300 167.815 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.615 3.300 161.215 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.315 3.300 157.915 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 162.915 3.300 164.515 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.400 3.300 245.000 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 236.800 3.300 238.400 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 240.100 3.300 241.700 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.500 3.300 235.100 211.800 ;
    END
  END vssa1
  PIN vssd1
    ANTENNADIFFAREA 15.428800 ;
    PORT
      LAYER met4 ;
        RECT 201.105 3.300 202.705 211.800 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER met4 ;
        RECT 213.440 3.300 215.040 211.800 ;
    END
  END vccd1
  OBS
      LAYER li1 ;
        RECT 144.605 64.060 276.725 133.815 ;
      LAYER met1 ;
        RECT 144.345 63.930 276.985 134.100 ;
      LAYER met2 ;
        RECT 7.745 165.585 515.545 166.965 ;
        RECT 7.745 142.040 515.825 165.585 ;
        RECT 7.465 65.210 515.825 142.040 ;
        RECT 7.465 64.435 203.500 65.210 ;
        RECT 7.465 0.000 199.300 64.435 ;
        RECT 200.140 0.000 203.500 64.435 ;
        RECT 204.340 0.000 215.915 65.210 ;
        RECT 216.755 0.000 515.825 65.210 ;
      LAYER met3 ;
        RECT 151.100 63.930 269.710 134.100 ;
  END
END sky130_ef_ip__xtal_osc_32k_DI
END LIBRARY

