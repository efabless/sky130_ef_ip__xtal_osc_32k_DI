magic
tech sky130A
magscale 1 2
timestamp 1527873355
<< checkpaint >>
rect 105 -1916 104553 44965
<< via1 >>
rect 29077 26665 29193 26781
rect 44245 26665 44361 26781
rect 39955 12831 40071 12947
<< metal2 >>
rect 1365 28664 1493 43705
rect 103165 33393 103293 43705
rect 44204 33173 103293 33393
rect 1365 28464 29235 28664
rect 29034 26781 29234 28464
rect 29034 26665 29077 26781
rect 29193 26665 29234 26781
rect 44204 26781 44404 33173
rect 29034 26620 29234 26665
rect 44204 26665 44245 26781
rect 44361 26665 44404 26781
rect 44204 26620 44404 26665
rect 39916 12947 40116 12986
rect 39916 12831 39955 12947
rect 40071 12831 40116 12947
rect 39916 0 40116 12831
rect 40756 0 40956 12863
rect 43239 0 43439 12863
rect 39916 -656 39972 0
rect 40756 -656 40812 0
rect 43239 -656 43295 0
<< via2 >>
rect 31269 26744 31325 26800
rect 31349 26744 31405 26800
rect 31429 26744 31485 26800
rect 31509 26744 31565 26800
rect 31935 26744 31991 26800
rect 32015 26744 32071 26800
rect 32095 26744 32151 26800
rect 32175 26744 32231 26800
rect 32594 26740 32650 26796
rect 32674 26740 32730 26796
rect 32754 26740 32810 26796
rect 32834 26740 32890 26796
rect 33257 26740 33313 26796
rect 33337 26740 33393 26796
rect 33417 26740 33473 26796
rect 33497 26740 33553 26796
rect 35398 26744 35454 26800
rect 35478 26744 35534 26800
rect 35558 26744 35614 26800
rect 35638 26744 35694 26800
rect 36064 26744 36120 26800
rect 36144 26744 36200 26800
rect 36224 26744 36280 26800
rect 36304 26744 36360 26800
rect 36723 26740 36779 26796
rect 36803 26740 36859 26796
rect 36883 26740 36939 26796
rect 36963 26740 37019 26796
rect 37386 26740 37442 26796
rect 37466 26740 37522 26796
rect 37546 26740 37602 26796
rect 37626 26740 37682 26796
rect 31269 26632 31325 26688
rect 31349 26632 31405 26688
rect 31429 26632 31485 26688
rect 31509 26632 31565 26688
rect 31935 26632 31991 26688
rect 32015 26632 32071 26688
rect 32095 26632 32151 26688
rect 32175 26632 32231 26688
rect 32594 26628 32650 26684
rect 32674 26628 32730 26684
rect 32754 26628 32810 26684
rect 32834 26628 32890 26684
rect 33257 26628 33313 26684
rect 33337 26628 33393 26684
rect 33417 26628 33473 26684
rect 33497 26628 33553 26684
rect 35398 26632 35454 26688
rect 35478 26632 35534 26688
rect 35558 26632 35614 26688
rect 35638 26632 35694 26688
rect 36064 26632 36120 26688
rect 36144 26632 36200 26688
rect 36224 26632 36280 26688
rect 36304 26632 36360 26688
rect 36723 26628 36779 26684
rect 36803 26628 36859 26684
rect 36883 26628 36939 26684
rect 36963 26628 37019 26684
rect 37386 26628 37442 26684
rect 37466 26628 37522 26684
rect 37546 26628 37602 26684
rect 37626 26628 37682 26684
rect 46706 26744 46762 26800
rect 46786 26744 46842 26800
rect 46866 26744 46922 26800
rect 46946 26744 47002 26800
rect 47372 26744 47428 26800
rect 47452 26744 47508 26800
rect 47532 26744 47588 26800
rect 47612 26744 47668 26800
rect 48031 26740 48087 26796
rect 48111 26740 48167 26796
rect 48191 26740 48247 26796
rect 48271 26740 48327 26796
rect 48694 26740 48750 26796
rect 48774 26740 48830 26796
rect 48854 26740 48910 26796
rect 48934 26740 48990 26796
rect 50835 26744 50891 26800
rect 50915 26744 50971 26800
rect 50995 26744 51051 26800
rect 51075 26744 51131 26800
rect 51501 26744 51557 26800
rect 51581 26744 51637 26800
rect 51661 26744 51717 26800
rect 51741 26744 51797 26800
rect 52160 26740 52216 26796
rect 52240 26740 52296 26796
rect 52320 26740 52376 26796
rect 52400 26740 52456 26796
rect 52823 26740 52879 26796
rect 52903 26740 52959 26796
rect 52983 26740 53039 26796
rect 53063 26740 53119 26796
rect 46706 26632 46762 26688
rect 46786 26632 46842 26688
rect 46866 26632 46922 26688
rect 46946 26632 47002 26688
rect 47372 26632 47428 26688
rect 47452 26632 47508 26688
rect 47532 26632 47588 26688
rect 47612 26632 47668 26688
rect 48031 26628 48087 26684
rect 48111 26628 48167 26684
rect 48191 26628 48247 26684
rect 48271 26628 48327 26684
rect 48694 26628 48750 26684
rect 48774 26628 48830 26684
rect 48854 26628 48910 26684
rect 48934 26628 48990 26684
rect 50835 26632 50891 26688
rect 50915 26632 50971 26688
rect 50995 26632 51051 26688
rect 51075 26632 51131 26688
rect 51501 26632 51557 26688
rect 51581 26632 51637 26688
rect 51661 26632 51717 26688
rect 51741 26632 51797 26688
rect 52160 26628 52216 26684
rect 52240 26628 52296 26684
rect 52320 26628 52376 26684
rect 52400 26628 52456 26684
rect 52823 26628 52879 26684
rect 52903 26628 52959 26684
rect 52983 26628 53039 26684
rect 53063 26628 53119 26684
rect 31269 26513 31325 26569
rect 31349 26513 31405 26569
rect 31429 26513 31485 26569
rect 31509 26513 31565 26569
rect 31935 26513 31991 26569
rect 32015 26513 32071 26569
rect 32095 26513 32151 26569
rect 32175 26513 32231 26569
rect 32594 26509 32650 26565
rect 32674 26509 32730 26565
rect 32754 26509 32810 26565
rect 32834 26509 32890 26565
rect 33257 26509 33313 26565
rect 33337 26509 33393 26565
rect 33417 26509 33473 26565
rect 33497 26509 33553 26565
rect 35398 26513 35454 26569
rect 35478 26513 35534 26569
rect 35558 26513 35614 26569
rect 35638 26513 35694 26569
rect 36064 26513 36120 26569
rect 36144 26513 36200 26569
rect 36224 26513 36280 26569
rect 36304 26513 36360 26569
rect 36723 26509 36779 26565
rect 36803 26509 36859 26565
rect 36883 26509 36939 26565
rect 36963 26509 37019 26565
rect 37386 26509 37442 26565
rect 37466 26509 37522 26565
rect 37546 26509 37602 26565
rect 37626 26509 37682 26565
rect 46706 26513 46762 26569
rect 46786 26513 46842 26569
rect 46866 26513 46922 26569
rect 46946 26513 47002 26569
rect 47372 26513 47428 26569
rect 47452 26513 47508 26569
rect 47532 26513 47588 26569
rect 47612 26513 47668 26569
rect 48031 26509 48087 26565
rect 48111 26509 48167 26565
rect 48191 26509 48247 26565
rect 48271 26509 48327 26565
rect 48694 26509 48750 26565
rect 48774 26509 48830 26565
rect 48854 26509 48910 26565
rect 48934 26509 48990 26565
rect 50835 26513 50891 26569
rect 50915 26513 50971 26569
rect 50995 26513 51051 26569
rect 51075 26513 51131 26569
rect 51501 26513 51557 26569
rect 51581 26513 51637 26569
rect 51661 26513 51717 26569
rect 51741 26513 51797 26569
rect 52160 26509 52216 26565
rect 52240 26509 52296 26565
rect 52320 26509 52376 26565
rect 52400 26509 52456 26565
rect 52823 26509 52879 26565
rect 52903 26509 52959 26565
rect 52983 26509 53039 26565
rect 53063 26509 53119 26565
rect 40319 13564 40375 13620
rect 40399 13564 40455 13620
rect 42794 13508 42850 13564
rect 42874 13508 42930 13564
rect 40319 13445 40375 13501
rect 40399 13445 40455 13501
rect 42794 13385 42850 13441
rect 42874 13385 42930 13441
rect 40319 13324 40375 13380
rect 40399 13324 40455 13380
rect 42794 13273 42850 13329
rect 42874 13273 42930 13329
rect 40319 13217 40375 13273
rect 40399 13217 40455 13273
rect 42794 13154 42850 13210
rect 42874 13154 42930 13210
rect 31269 13052 31325 13108
rect 31349 13052 31405 13108
rect 31429 13052 31485 13108
rect 31509 13052 31565 13108
rect 31935 13052 31991 13108
rect 32015 13052 32071 13108
rect 32095 13052 32151 13108
rect 32175 13052 32231 13108
rect 32594 13048 32650 13104
rect 32674 13048 32730 13104
rect 32754 13048 32810 13104
rect 32834 13048 32890 13104
rect 33257 13048 33313 13104
rect 33337 13048 33393 13104
rect 33417 13048 33473 13104
rect 33497 13048 33553 13104
rect 35398 13052 35454 13108
rect 35478 13052 35534 13108
rect 35558 13052 35614 13108
rect 35638 13052 35694 13108
rect 36064 13052 36120 13108
rect 36144 13052 36200 13108
rect 36224 13052 36280 13108
rect 36304 13052 36360 13108
rect 36723 13048 36779 13104
rect 36803 13048 36859 13104
rect 36883 13048 36939 13104
rect 36963 13048 37019 13104
rect 37386 13048 37442 13104
rect 37466 13048 37522 13104
rect 37546 13048 37602 13104
rect 37626 13048 37682 13104
rect 40319 13091 40375 13147
rect 40399 13091 40455 13147
rect 31269 12940 31325 12996
rect 31349 12940 31405 12996
rect 31429 12940 31485 12996
rect 31509 12940 31565 12996
rect 31935 12940 31991 12996
rect 32015 12940 32071 12996
rect 32095 12940 32151 12996
rect 32175 12940 32231 12996
rect 32594 12936 32650 12992
rect 32674 12936 32730 12992
rect 32754 12936 32810 12992
rect 32834 12936 32890 12992
rect 33257 12936 33313 12992
rect 33337 12936 33393 12992
rect 33417 12936 33473 12992
rect 33497 12936 33553 12992
rect 35398 12940 35454 12996
rect 35478 12940 35534 12996
rect 35558 12940 35614 12996
rect 35638 12940 35694 12996
rect 36064 12940 36120 12996
rect 36144 12940 36200 12996
rect 36224 12940 36280 12996
rect 36304 12940 36360 12996
rect 36723 12936 36779 12992
rect 36803 12936 36859 12992
rect 36883 12936 36939 12992
rect 36963 12936 37019 12992
rect 37386 12936 37442 12992
rect 37466 12936 37522 12992
rect 37546 12936 37602 12992
rect 37626 12936 37682 12992
rect 40319 12979 40375 13035
rect 40399 12979 40455 13035
rect 42794 13030 42850 13086
rect 42874 13030 42930 13086
rect 46706 13052 46762 13108
rect 46786 13052 46842 13108
rect 46866 13052 46922 13108
rect 46946 13052 47002 13108
rect 47372 13052 47428 13108
rect 47452 13052 47508 13108
rect 47532 13052 47588 13108
rect 47612 13052 47668 13108
rect 48031 13048 48087 13104
rect 48111 13048 48167 13104
rect 48191 13048 48247 13104
rect 48271 13048 48327 13104
rect 48694 13048 48750 13104
rect 48774 13048 48830 13104
rect 48854 13048 48910 13104
rect 48934 13048 48990 13104
rect 50835 13052 50891 13108
rect 50915 13052 50971 13108
rect 50995 13052 51051 13108
rect 51075 13052 51131 13108
rect 51501 13052 51557 13108
rect 51581 13052 51637 13108
rect 51661 13052 51717 13108
rect 51741 13052 51797 13108
rect 52160 13048 52216 13104
rect 52240 13048 52296 13104
rect 52320 13048 52376 13104
rect 52400 13048 52456 13104
rect 52823 13048 52879 13104
rect 52903 13048 52959 13104
rect 52983 13048 53039 13104
rect 53063 13048 53119 13104
rect 31269 12821 31325 12877
rect 31349 12821 31405 12877
rect 31429 12821 31485 12877
rect 31509 12821 31565 12877
rect 31935 12821 31991 12877
rect 32015 12821 32071 12877
rect 32095 12821 32151 12877
rect 32175 12821 32231 12877
rect 32594 12817 32650 12873
rect 32674 12817 32730 12873
rect 32754 12817 32810 12873
rect 32834 12817 32890 12873
rect 33257 12817 33313 12873
rect 33337 12817 33393 12873
rect 33417 12817 33473 12873
rect 33497 12817 33553 12873
rect 35398 12821 35454 12877
rect 35478 12821 35534 12877
rect 35558 12821 35614 12877
rect 35638 12821 35694 12877
rect 36064 12821 36120 12877
rect 36144 12821 36200 12877
rect 36224 12821 36280 12877
rect 36304 12821 36360 12877
rect 36723 12817 36779 12873
rect 36803 12817 36859 12873
rect 36883 12817 36939 12873
rect 36963 12817 37019 12873
rect 37386 12817 37442 12873
rect 37466 12817 37522 12873
rect 37546 12817 37602 12873
rect 37626 12817 37682 12873
rect 42794 12923 42850 12979
rect 42874 12923 42930 12979
rect 46706 12940 46762 12996
rect 46786 12940 46842 12996
rect 46866 12940 46922 12996
rect 46946 12940 47002 12996
rect 47372 12940 47428 12996
rect 47452 12940 47508 12996
rect 47532 12940 47588 12996
rect 47612 12940 47668 12996
rect 48031 12936 48087 12992
rect 48111 12936 48167 12992
rect 48191 12936 48247 12992
rect 48271 12936 48327 12992
rect 48694 12936 48750 12992
rect 48774 12936 48830 12992
rect 48854 12936 48910 12992
rect 48934 12936 48990 12992
rect 50835 12940 50891 12996
rect 50915 12940 50971 12996
rect 50995 12940 51051 12996
rect 51075 12940 51131 12996
rect 51501 12940 51557 12996
rect 51581 12940 51637 12996
rect 51661 12940 51717 12996
rect 51741 12940 51797 12996
rect 52160 12936 52216 12992
rect 52240 12936 52296 12992
rect 52320 12936 52376 12992
rect 52400 12936 52456 12992
rect 52823 12936 52879 12992
rect 52903 12936 52959 12992
rect 52983 12936 53039 12992
rect 53063 12936 53119 12992
rect 40319 12860 40375 12916
rect 40399 12860 40455 12916
rect 46706 12821 46762 12877
rect 46786 12821 46842 12877
rect 46866 12821 46922 12877
rect 46946 12821 47002 12877
rect 47372 12821 47428 12877
rect 47452 12821 47508 12877
rect 47532 12821 47588 12877
rect 47612 12821 47668 12877
rect 48031 12817 48087 12873
rect 48111 12817 48167 12873
rect 48191 12817 48247 12873
rect 48271 12817 48327 12873
rect 48694 12817 48750 12873
rect 48774 12817 48830 12873
rect 48854 12817 48910 12873
rect 48934 12817 48990 12873
rect 50835 12821 50891 12877
rect 50915 12821 50971 12877
rect 50995 12821 51051 12877
rect 51075 12821 51131 12877
rect 51501 12821 51557 12877
rect 51581 12821 51637 12877
rect 51661 12821 51717 12877
rect 51741 12821 51797 12877
rect 52160 12817 52216 12873
rect 52240 12817 52296 12873
rect 52320 12817 52376 12873
rect 52400 12817 52456 12873
rect 52823 12817 52879 12873
rect 52903 12817 52959 12873
rect 52983 12817 53039 12873
rect 53063 12817 53119 12873
<< metal3 >>
rect 30220 26804 34220 26820
rect 30220 26740 31265 26804
rect 31329 26740 31345 26804
rect 31409 26740 31425 26804
rect 31489 26740 31505 26804
rect 31569 26740 31931 26804
rect 31995 26740 32011 26804
rect 32075 26740 32091 26804
rect 32155 26740 32171 26804
rect 32235 26800 34220 26804
rect 32235 26740 32590 26800
rect 30220 26736 32590 26740
rect 32654 26736 32670 26800
rect 32734 26736 32750 26800
rect 32814 26736 32830 26800
rect 32894 26736 33253 26800
rect 33317 26736 33333 26800
rect 33397 26736 33413 26800
rect 33477 26736 33493 26800
rect 33557 26736 34220 26800
rect 30220 26692 34220 26736
rect 30220 26628 31265 26692
rect 31329 26628 31345 26692
rect 31409 26628 31425 26692
rect 31489 26628 31505 26692
rect 31569 26628 31931 26692
rect 31995 26628 32011 26692
rect 32075 26628 32091 26692
rect 32155 26628 32171 26692
rect 32235 26688 34220 26692
rect 32235 26628 32590 26688
rect 30220 26624 32590 26628
rect 32654 26624 32670 26688
rect 32734 26624 32750 26688
rect 32814 26624 32830 26688
rect 32894 26624 33253 26688
rect 33317 26624 33333 26688
rect 33397 26624 33413 26688
rect 33477 26624 33493 26688
rect 33557 26624 34220 26688
rect 30220 26573 34220 26624
rect 30220 26509 31265 26573
rect 31329 26509 31345 26573
rect 31409 26509 31425 26573
rect 31489 26509 31505 26573
rect 31569 26509 31931 26573
rect 31995 26509 32011 26573
rect 32075 26509 32091 26573
rect 32155 26509 32171 26573
rect 32235 26569 34220 26573
rect 32235 26509 32590 26569
rect 30220 26505 32590 26509
rect 32654 26505 32670 26569
rect 32734 26505 32750 26569
rect 32814 26505 32830 26569
rect 32894 26505 33253 26569
rect 33317 26505 33333 26569
rect 33397 26505 33413 26569
rect 33477 26505 33493 26569
rect 33557 26505 34220 26569
rect 30220 26478 34220 26505
rect 34505 26804 38505 26820
rect 34505 26740 35394 26804
rect 35458 26740 35474 26804
rect 35538 26740 35554 26804
rect 35618 26740 35634 26804
rect 35698 26740 36060 26804
rect 36124 26740 36140 26804
rect 36204 26740 36220 26804
rect 36284 26740 36300 26804
rect 36364 26800 38505 26804
rect 36364 26740 36719 26800
rect 34505 26736 36719 26740
rect 36783 26736 36799 26800
rect 36863 26736 36879 26800
rect 36943 26736 36959 26800
rect 37023 26736 37382 26800
rect 37446 26736 37462 26800
rect 37526 26736 37542 26800
rect 37606 26736 37622 26800
rect 37686 26736 38505 26800
rect 34505 26692 38505 26736
rect 34505 26628 35394 26692
rect 35458 26628 35474 26692
rect 35538 26628 35554 26692
rect 35618 26628 35634 26692
rect 35698 26628 36060 26692
rect 36124 26628 36140 26692
rect 36204 26628 36220 26692
rect 36284 26628 36300 26692
rect 36364 26688 38505 26692
rect 36364 26628 36719 26688
rect 34505 26624 36719 26628
rect 36783 26624 36799 26688
rect 36863 26624 36879 26688
rect 36943 26624 36959 26688
rect 37023 26624 37382 26688
rect 37446 26624 37462 26688
rect 37526 26624 37542 26688
rect 37606 26624 37622 26688
rect 37686 26624 38505 26688
rect 34505 26573 38505 26624
rect 34505 26509 35394 26573
rect 35458 26509 35474 26573
rect 35538 26509 35554 26573
rect 35618 26509 35634 26573
rect 35698 26509 36060 26573
rect 36124 26509 36140 26573
rect 36204 26509 36220 26573
rect 36284 26509 36300 26573
rect 36364 26569 38505 26573
rect 36364 26509 36719 26569
rect 34505 26505 36719 26509
rect 36783 26505 36799 26569
rect 36863 26505 36879 26569
rect 36943 26505 36959 26569
rect 37023 26505 37382 26569
rect 37446 26505 37462 26569
rect 37526 26505 37542 26569
rect 37606 26505 37622 26569
rect 37686 26505 38505 26569
rect 34505 26478 38505 26505
rect 45657 26804 49657 26820
rect 45657 26740 46702 26804
rect 46766 26740 46782 26804
rect 46846 26740 46862 26804
rect 46926 26740 46942 26804
rect 47006 26740 47368 26804
rect 47432 26740 47448 26804
rect 47512 26740 47528 26804
rect 47592 26740 47608 26804
rect 47672 26800 49657 26804
rect 47672 26740 48027 26800
rect 45657 26736 48027 26740
rect 48091 26736 48107 26800
rect 48171 26736 48187 26800
rect 48251 26736 48267 26800
rect 48331 26736 48690 26800
rect 48754 26736 48770 26800
rect 48834 26736 48850 26800
rect 48914 26736 48930 26800
rect 48994 26736 49657 26800
rect 45657 26692 49657 26736
rect 45657 26628 46702 26692
rect 46766 26628 46782 26692
rect 46846 26628 46862 26692
rect 46926 26628 46942 26692
rect 47006 26628 47368 26692
rect 47432 26628 47448 26692
rect 47512 26628 47528 26692
rect 47592 26628 47608 26692
rect 47672 26688 49657 26692
rect 47672 26628 48027 26688
rect 45657 26624 48027 26628
rect 48091 26624 48107 26688
rect 48171 26624 48187 26688
rect 48251 26624 48267 26688
rect 48331 26624 48690 26688
rect 48754 26624 48770 26688
rect 48834 26624 48850 26688
rect 48914 26624 48930 26688
rect 48994 26624 49657 26688
rect 45657 26573 49657 26624
rect 45657 26509 46702 26573
rect 46766 26509 46782 26573
rect 46846 26509 46862 26573
rect 46926 26509 46942 26573
rect 47006 26509 47368 26573
rect 47432 26509 47448 26573
rect 47512 26509 47528 26573
rect 47592 26509 47608 26573
rect 47672 26569 49657 26573
rect 47672 26509 48027 26569
rect 45657 26505 48027 26509
rect 48091 26505 48107 26569
rect 48171 26505 48187 26569
rect 48251 26505 48267 26569
rect 48331 26505 48690 26569
rect 48754 26505 48770 26569
rect 48834 26505 48850 26569
rect 48914 26505 48930 26569
rect 48994 26505 49657 26569
rect 45657 26478 49657 26505
rect 49942 26804 53942 26820
rect 49942 26740 50831 26804
rect 50895 26740 50911 26804
rect 50975 26740 50991 26804
rect 51055 26740 51071 26804
rect 51135 26740 51497 26804
rect 51561 26740 51577 26804
rect 51641 26740 51657 26804
rect 51721 26740 51737 26804
rect 51801 26800 53942 26804
rect 51801 26740 52156 26800
rect 49942 26736 52156 26740
rect 52220 26736 52236 26800
rect 52300 26736 52316 26800
rect 52380 26736 52396 26800
rect 52460 26736 52819 26800
rect 52883 26736 52899 26800
rect 52963 26736 52979 26800
rect 53043 26736 53059 26800
rect 53123 26736 53942 26800
rect 49942 26692 53942 26736
rect 49942 26628 50831 26692
rect 50895 26628 50911 26692
rect 50975 26628 50991 26692
rect 51055 26628 51071 26692
rect 51135 26628 51497 26692
rect 51561 26628 51577 26692
rect 51641 26628 51657 26692
rect 51721 26628 51737 26692
rect 51801 26688 53942 26692
rect 51801 26628 52156 26688
rect 49942 26624 52156 26628
rect 52220 26624 52236 26688
rect 52300 26624 52316 26688
rect 52380 26624 52396 26688
rect 52460 26624 52819 26688
rect 52883 26624 52899 26688
rect 52963 26624 52979 26688
rect 53043 26624 53059 26688
rect 53123 26624 53942 26688
rect 49942 26573 53942 26624
rect 49942 26509 50831 26573
rect 50895 26509 50911 26573
rect 50975 26509 50991 26573
rect 51055 26509 51071 26573
rect 51135 26509 51497 26573
rect 51561 26509 51577 26573
rect 51641 26509 51657 26573
rect 51721 26509 51737 26573
rect 51801 26569 53942 26573
rect 51801 26509 52156 26569
rect 49942 26505 52156 26509
rect 52220 26505 52236 26569
rect 52300 26505 52316 26569
rect 52380 26505 52396 26569
rect 52460 26505 52819 26569
rect 52883 26505 52899 26569
rect 52963 26505 52979 26569
rect 53043 26505 53059 26569
rect 53123 26505 53942 26569
rect 49942 26478 53942 26505
rect 40279 13624 40479 13718
rect 40279 13560 40315 13624
rect 40379 13560 40395 13624
rect 40459 13560 40479 13624
rect 40279 13505 40479 13560
rect 40279 13441 40315 13505
rect 40379 13441 40395 13505
rect 40459 13441 40479 13505
rect 40279 13384 40479 13441
rect 40279 13320 40315 13384
rect 40379 13320 40395 13384
rect 40459 13320 40479 13384
rect 40279 13277 40479 13320
rect 40279 13213 40315 13277
rect 40379 13213 40395 13277
rect 40459 13213 40479 13277
rect 40279 13151 40479 13213
rect 30220 13112 34220 13128
rect 30220 13048 31265 13112
rect 31329 13048 31345 13112
rect 31409 13048 31425 13112
rect 31489 13048 31505 13112
rect 31569 13048 31931 13112
rect 31995 13048 32011 13112
rect 32075 13048 32091 13112
rect 32155 13048 32171 13112
rect 32235 13108 34220 13112
rect 32235 13048 32590 13108
rect 30220 13044 32590 13048
rect 32654 13044 32670 13108
rect 32734 13044 32750 13108
rect 32814 13044 32830 13108
rect 32894 13044 33253 13108
rect 33317 13044 33333 13108
rect 33397 13044 33413 13108
rect 33477 13044 33493 13108
rect 33557 13044 34220 13108
rect 30220 13000 34220 13044
rect 30220 12936 31265 13000
rect 31329 12936 31345 13000
rect 31409 12936 31425 13000
rect 31489 12936 31505 13000
rect 31569 12936 31931 13000
rect 31995 12936 32011 13000
rect 32075 12936 32091 13000
rect 32155 12936 32171 13000
rect 32235 12996 34220 13000
rect 32235 12936 32590 12996
rect 30220 12932 32590 12936
rect 32654 12932 32670 12996
rect 32734 12932 32750 12996
rect 32814 12932 32830 12996
rect 32894 12932 33253 12996
rect 33317 12932 33333 12996
rect 33397 12932 33413 12996
rect 33477 12932 33493 12996
rect 33557 12932 34220 12996
rect 30220 12881 34220 12932
rect 30220 12817 31265 12881
rect 31329 12817 31345 12881
rect 31409 12817 31425 12881
rect 31489 12817 31505 12881
rect 31569 12817 31931 12881
rect 31995 12817 32011 12881
rect 32075 12817 32091 12881
rect 32155 12817 32171 12881
rect 32235 12877 34220 12881
rect 32235 12817 32590 12877
rect 30220 12813 32590 12817
rect 32654 12813 32670 12877
rect 32734 12813 32750 12877
rect 32814 12813 32830 12877
rect 32894 12813 33253 12877
rect 33317 12813 33333 12877
rect 33397 12813 33413 12877
rect 33477 12813 33493 12877
rect 33557 12813 34220 12877
rect 30220 12786 34220 12813
rect 34505 13112 38505 13128
rect 34505 13048 35394 13112
rect 35458 13048 35474 13112
rect 35538 13048 35554 13112
rect 35618 13048 35634 13112
rect 35698 13048 36060 13112
rect 36124 13048 36140 13112
rect 36204 13048 36220 13112
rect 36284 13048 36300 13112
rect 36364 13108 38505 13112
rect 36364 13048 36719 13108
rect 34505 13044 36719 13048
rect 36783 13044 36799 13108
rect 36863 13044 36879 13108
rect 36943 13044 36959 13108
rect 37023 13044 37382 13108
rect 37446 13044 37462 13108
rect 37526 13044 37542 13108
rect 37606 13044 37622 13108
rect 37686 13044 38505 13108
rect 34505 13000 38505 13044
rect 34505 12936 35394 13000
rect 35458 12936 35474 13000
rect 35538 12936 35554 13000
rect 35618 12936 35634 13000
rect 35698 12936 36060 13000
rect 36124 12936 36140 13000
rect 36204 12936 36220 13000
rect 36284 12936 36300 13000
rect 36364 12996 38505 13000
rect 36364 12936 36719 12996
rect 34505 12932 36719 12936
rect 36783 12932 36799 12996
rect 36863 12932 36879 12996
rect 36943 12932 36959 12996
rect 37023 12932 37382 12996
rect 37446 12932 37462 12996
rect 37526 12932 37542 12996
rect 37606 12932 37622 12996
rect 37686 12932 38505 12996
rect 34505 12881 38505 12932
rect 34505 12817 35394 12881
rect 35458 12817 35474 12881
rect 35538 12817 35554 12881
rect 35618 12817 35634 12881
rect 35698 12817 36060 12881
rect 36124 12817 36140 12881
rect 36204 12817 36220 12881
rect 36284 12817 36300 12881
rect 36364 12877 38505 12881
rect 36364 12817 36719 12877
rect 34505 12813 36719 12817
rect 36783 12813 36799 12877
rect 36863 12813 36879 12877
rect 36943 12813 36959 12877
rect 37023 12813 37382 12877
rect 37446 12813 37462 12877
rect 37526 12813 37542 12877
rect 37606 12813 37622 12877
rect 37686 12813 38505 12877
rect 34505 12786 38505 12813
rect 40279 13087 40315 13151
rect 40379 13087 40395 13151
rect 40459 13087 40479 13151
rect 40279 13039 40479 13087
rect 40279 12975 40315 13039
rect 40379 12975 40395 13039
rect 40459 12975 40479 13039
rect 40279 12920 40479 12975
rect 40279 12856 40315 12920
rect 40379 12856 40395 12920
rect 40459 12856 40479 12920
rect 40279 12786 40479 12856
rect 42754 13568 42954 13575
rect 42754 13504 42790 13568
rect 42854 13504 42870 13568
rect 42934 13504 42954 13568
rect 42754 13445 42954 13504
rect 42754 13381 42790 13445
rect 42854 13381 42870 13445
rect 42934 13381 42954 13445
rect 42754 13333 42954 13381
rect 42754 13269 42790 13333
rect 42854 13269 42870 13333
rect 42934 13269 42954 13333
rect 42754 13214 42954 13269
rect 42754 13150 42790 13214
rect 42854 13150 42870 13214
rect 42934 13150 42954 13214
rect 42754 13090 42954 13150
rect 42754 13026 42790 13090
rect 42854 13026 42870 13090
rect 42934 13026 42954 13090
rect 42754 12983 42954 13026
rect 42754 12919 42790 12983
rect 42854 12919 42870 12983
rect 42934 12919 42954 12983
rect 42754 12786 42954 12919
rect 45657 13112 49657 13128
rect 45657 13048 46702 13112
rect 46766 13048 46782 13112
rect 46846 13048 46862 13112
rect 46926 13048 46942 13112
rect 47006 13048 47368 13112
rect 47432 13048 47448 13112
rect 47512 13048 47528 13112
rect 47592 13048 47608 13112
rect 47672 13108 49657 13112
rect 47672 13048 48027 13108
rect 45657 13044 48027 13048
rect 48091 13044 48107 13108
rect 48171 13044 48187 13108
rect 48251 13044 48267 13108
rect 48331 13044 48690 13108
rect 48754 13044 48770 13108
rect 48834 13044 48850 13108
rect 48914 13044 48930 13108
rect 48994 13044 49657 13108
rect 45657 13000 49657 13044
rect 45657 12936 46702 13000
rect 46766 12936 46782 13000
rect 46846 12936 46862 13000
rect 46926 12936 46942 13000
rect 47006 12936 47368 13000
rect 47432 12936 47448 13000
rect 47512 12936 47528 13000
rect 47592 12936 47608 13000
rect 47672 12996 49657 13000
rect 47672 12936 48027 12996
rect 45657 12932 48027 12936
rect 48091 12932 48107 12996
rect 48171 12932 48187 12996
rect 48251 12932 48267 12996
rect 48331 12932 48690 12996
rect 48754 12932 48770 12996
rect 48834 12932 48850 12996
rect 48914 12932 48930 12996
rect 48994 12932 49657 12996
rect 45657 12881 49657 12932
rect 45657 12817 46702 12881
rect 46766 12817 46782 12881
rect 46846 12817 46862 12881
rect 46926 12817 46942 12881
rect 47006 12817 47368 12881
rect 47432 12817 47448 12881
rect 47512 12817 47528 12881
rect 47592 12817 47608 12881
rect 47672 12877 49657 12881
rect 47672 12817 48027 12877
rect 45657 12813 48027 12817
rect 48091 12813 48107 12877
rect 48171 12813 48187 12877
rect 48251 12813 48267 12877
rect 48331 12813 48690 12877
rect 48754 12813 48770 12877
rect 48834 12813 48850 12877
rect 48914 12813 48930 12877
rect 48994 12813 49657 12877
rect 45657 12786 49657 12813
rect 49942 13112 53942 13128
rect 49942 13048 50831 13112
rect 50895 13048 50911 13112
rect 50975 13048 50991 13112
rect 51055 13048 51071 13112
rect 51135 13048 51497 13112
rect 51561 13048 51577 13112
rect 51641 13048 51657 13112
rect 51721 13048 51737 13112
rect 51801 13108 53942 13112
rect 51801 13048 52156 13108
rect 49942 13044 52156 13048
rect 52220 13044 52236 13108
rect 52300 13044 52316 13108
rect 52380 13044 52396 13108
rect 52460 13044 52819 13108
rect 52883 13044 52899 13108
rect 52963 13044 52979 13108
rect 53043 13044 53059 13108
rect 53123 13044 53942 13108
rect 49942 13000 53942 13044
rect 49942 12936 50831 13000
rect 50895 12936 50911 13000
rect 50975 12936 50991 13000
rect 51055 12936 51071 13000
rect 51135 12936 51497 13000
rect 51561 12936 51577 13000
rect 51641 12936 51657 13000
rect 51721 12936 51737 13000
rect 51801 12996 53942 13000
rect 51801 12936 52156 12996
rect 49942 12932 52156 12936
rect 52220 12932 52236 12996
rect 52300 12932 52316 12996
rect 52380 12932 52396 12996
rect 52460 12932 52819 12996
rect 52883 12932 52899 12996
rect 52963 12932 52979 12996
rect 53043 12932 53059 12996
rect 53123 12932 53942 12996
rect 49942 12881 53942 12932
rect 49942 12817 50831 12881
rect 50895 12817 50911 12881
rect 50975 12817 50991 12881
rect 51055 12817 51071 12881
rect 51135 12817 51497 12881
rect 51561 12817 51577 12881
rect 51641 12817 51657 12881
rect 51721 12817 51737 12881
rect 51801 12877 53942 12881
rect 51801 12817 52156 12877
rect 49942 12813 52156 12817
rect 52220 12813 52236 12877
rect 52300 12813 52316 12877
rect 52380 12813 52396 12877
rect 52460 12813 52819 12877
rect 52883 12813 52899 12877
rect 52963 12813 52979 12877
rect 53043 12813 53059 12877
rect 53123 12813 53942 12877
rect 49942 12786 53942 12813
<< via3 >>
rect 31265 26800 31329 26804
rect 31265 26744 31269 26800
rect 31269 26744 31325 26800
rect 31325 26744 31329 26800
rect 31265 26740 31329 26744
rect 31345 26800 31409 26804
rect 31345 26744 31349 26800
rect 31349 26744 31405 26800
rect 31405 26744 31409 26800
rect 31345 26740 31409 26744
rect 31425 26800 31489 26804
rect 31425 26744 31429 26800
rect 31429 26744 31485 26800
rect 31485 26744 31489 26800
rect 31425 26740 31489 26744
rect 31505 26800 31569 26804
rect 31505 26744 31509 26800
rect 31509 26744 31565 26800
rect 31565 26744 31569 26800
rect 31505 26740 31569 26744
rect 31931 26800 31995 26804
rect 31931 26744 31935 26800
rect 31935 26744 31991 26800
rect 31991 26744 31995 26800
rect 31931 26740 31995 26744
rect 32011 26800 32075 26804
rect 32011 26744 32015 26800
rect 32015 26744 32071 26800
rect 32071 26744 32075 26800
rect 32011 26740 32075 26744
rect 32091 26800 32155 26804
rect 32091 26744 32095 26800
rect 32095 26744 32151 26800
rect 32151 26744 32155 26800
rect 32091 26740 32155 26744
rect 32171 26800 32235 26804
rect 32171 26744 32175 26800
rect 32175 26744 32231 26800
rect 32231 26744 32235 26800
rect 32171 26740 32235 26744
rect 32590 26796 32654 26800
rect 32590 26740 32594 26796
rect 32594 26740 32650 26796
rect 32650 26740 32654 26796
rect 32590 26736 32654 26740
rect 32670 26796 32734 26800
rect 32670 26740 32674 26796
rect 32674 26740 32730 26796
rect 32730 26740 32734 26796
rect 32670 26736 32734 26740
rect 32750 26796 32814 26800
rect 32750 26740 32754 26796
rect 32754 26740 32810 26796
rect 32810 26740 32814 26796
rect 32750 26736 32814 26740
rect 32830 26796 32894 26800
rect 32830 26740 32834 26796
rect 32834 26740 32890 26796
rect 32890 26740 32894 26796
rect 32830 26736 32894 26740
rect 33253 26796 33317 26800
rect 33253 26740 33257 26796
rect 33257 26740 33313 26796
rect 33313 26740 33317 26796
rect 33253 26736 33317 26740
rect 33333 26796 33397 26800
rect 33333 26740 33337 26796
rect 33337 26740 33393 26796
rect 33393 26740 33397 26796
rect 33333 26736 33397 26740
rect 33413 26796 33477 26800
rect 33413 26740 33417 26796
rect 33417 26740 33473 26796
rect 33473 26740 33477 26796
rect 33413 26736 33477 26740
rect 33493 26796 33557 26800
rect 33493 26740 33497 26796
rect 33497 26740 33553 26796
rect 33553 26740 33557 26796
rect 33493 26736 33557 26740
rect 31265 26688 31329 26692
rect 31265 26632 31269 26688
rect 31269 26632 31325 26688
rect 31325 26632 31329 26688
rect 31265 26628 31329 26632
rect 31345 26688 31409 26692
rect 31345 26632 31349 26688
rect 31349 26632 31405 26688
rect 31405 26632 31409 26688
rect 31345 26628 31409 26632
rect 31425 26688 31489 26692
rect 31425 26632 31429 26688
rect 31429 26632 31485 26688
rect 31485 26632 31489 26688
rect 31425 26628 31489 26632
rect 31505 26688 31569 26692
rect 31505 26632 31509 26688
rect 31509 26632 31565 26688
rect 31565 26632 31569 26688
rect 31505 26628 31569 26632
rect 31931 26688 31995 26692
rect 31931 26632 31935 26688
rect 31935 26632 31991 26688
rect 31991 26632 31995 26688
rect 31931 26628 31995 26632
rect 32011 26688 32075 26692
rect 32011 26632 32015 26688
rect 32015 26632 32071 26688
rect 32071 26632 32075 26688
rect 32011 26628 32075 26632
rect 32091 26688 32155 26692
rect 32091 26632 32095 26688
rect 32095 26632 32151 26688
rect 32151 26632 32155 26688
rect 32091 26628 32155 26632
rect 32171 26688 32235 26692
rect 32171 26632 32175 26688
rect 32175 26632 32231 26688
rect 32231 26632 32235 26688
rect 32171 26628 32235 26632
rect 32590 26684 32654 26688
rect 32590 26628 32594 26684
rect 32594 26628 32650 26684
rect 32650 26628 32654 26684
rect 32590 26624 32654 26628
rect 32670 26684 32734 26688
rect 32670 26628 32674 26684
rect 32674 26628 32730 26684
rect 32730 26628 32734 26684
rect 32670 26624 32734 26628
rect 32750 26684 32814 26688
rect 32750 26628 32754 26684
rect 32754 26628 32810 26684
rect 32810 26628 32814 26684
rect 32750 26624 32814 26628
rect 32830 26684 32894 26688
rect 32830 26628 32834 26684
rect 32834 26628 32890 26684
rect 32890 26628 32894 26684
rect 32830 26624 32894 26628
rect 33253 26684 33317 26688
rect 33253 26628 33257 26684
rect 33257 26628 33313 26684
rect 33313 26628 33317 26684
rect 33253 26624 33317 26628
rect 33333 26684 33397 26688
rect 33333 26628 33337 26684
rect 33337 26628 33393 26684
rect 33393 26628 33397 26684
rect 33333 26624 33397 26628
rect 33413 26684 33477 26688
rect 33413 26628 33417 26684
rect 33417 26628 33473 26684
rect 33473 26628 33477 26684
rect 33413 26624 33477 26628
rect 33493 26684 33557 26688
rect 33493 26628 33497 26684
rect 33497 26628 33553 26684
rect 33553 26628 33557 26684
rect 33493 26624 33557 26628
rect 31265 26569 31329 26573
rect 31265 26513 31269 26569
rect 31269 26513 31325 26569
rect 31325 26513 31329 26569
rect 31265 26509 31329 26513
rect 31345 26569 31409 26573
rect 31345 26513 31349 26569
rect 31349 26513 31405 26569
rect 31405 26513 31409 26569
rect 31345 26509 31409 26513
rect 31425 26569 31489 26573
rect 31425 26513 31429 26569
rect 31429 26513 31485 26569
rect 31485 26513 31489 26569
rect 31425 26509 31489 26513
rect 31505 26569 31569 26573
rect 31505 26513 31509 26569
rect 31509 26513 31565 26569
rect 31565 26513 31569 26569
rect 31505 26509 31569 26513
rect 31931 26569 31995 26573
rect 31931 26513 31935 26569
rect 31935 26513 31991 26569
rect 31991 26513 31995 26569
rect 31931 26509 31995 26513
rect 32011 26569 32075 26573
rect 32011 26513 32015 26569
rect 32015 26513 32071 26569
rect 32071 26513 32075 26569
rect 32011 26509 32075 26513
rect 32091 26569 32155 26573
rect 32091 26513 32095 26569
rect 32095 26513 32151 26569
rect 32151 26513 32155 26569
rect 32091 26509 32155 26513
rect 32171 26569 32235 26573
rect 32171 26513 32175 26569
rect 32175 26513 32231 26569
rect 32231 26513 32235 26569
rect 32171 26509 32235 26513
rect 32590 26565 32654 26569
rect 32590 26509 32594 26565
rect 32594 26509 32650 26565
rect 32650 26509 32654 26565
rect 32590 26505 32654 26509
rect 32670 26565 32734 26569
rect 32670 26509 32674 26565
rect 32674 26509 32730 26565
rect 32730 26509 32734 26565
rect 32670 26505 32734 26509
rect 32750 26565 32814 26569
rect 32750 26509 32754 26565
rect 32754 26509 32810 26565
rect 32810 26509 32814 26565
rect 32750 26505 32814 26509
rect 32830 26565 32894 26569
rect 32830 26509 32834 26565
rect 32834 26509 32890 26565
rect 32890 26509 32894 26565
rect 32830 26505 32894 26509
rect 33253 26565 33317 26569
rect 33253 26509 33257 26565
rect 33257 26509 33313 26565
rect 33313 26509 33317 26565
rect 33253 26505 33317 26509
rect 33333 26565 33397 26569
rect 33333 26509 33337 26565
rect 33337 26509 33393 26565
rect 33393 26509 33397 26565
rect 33333 26505 33397 26509
rect 33413 26565 33477 26569
rect 33413 26509 33417 26565
rect 33417 26509 33473 26565
rect 33473 26509 33477 26565
rect 33413 26505 33477 26509
rect 33493 26565 33557 26569
rect 33493 26509 33497 26565
rect 33497 26509 33553 26565
rect 33553 26509 33557 26565
rect 33493 26505 33557 26509
rect 35394 26800 35458 26804
rect 35394 26744 35398 26800
rect 35398 26744 35454 26800
rect 35454 26744 35458 26800
rect 35394 26740 35458 26744
rect 35474 26800 35538 26804
rect 35474 26744 35478 26800
rect 35478 26744 35534 26800
rect 35534 26744 35538 26800
rect 35474 26740 35538 26744
rect 35554 26800 35618 26804
rect 35554 26744 35558 26800
rect 35558 26744 35614 26800
rect 35614 26744 35618 26800
rect 35554 26740 35618 26744
rect 35634 26800 35698 26804
rect 35634 26744 35638 26800
rect 35638 26744 35694 26800
rect 35694 26744 35698 26800
rect 35634 26740 35698 26744
rect 36060 26800 36124 26804
rect 36060 26744 36064 26800
rect 36064 26744 36120 26800
rect 36120 26744 36124 26800
rect 36060 26740 36124 26744
rect 36140 26800 36204 26804
rect 36140 26744 36144 26800
rect 36144 26744 36200 26800
rect 36200 26744 36204 26800
rect 36140 26740 36204 26744
rect 36220 26800 36284 26804
rect 36220 26744 36224 26800
rect 36224 26744 36280 26800
rect 36280 26744 36284 26800
rect 36220 26740 36284 26744
rect 36300 26800 36364 26804
rect 36300 26744 36304 26800
rect 36304 26744 36360 26800
rect 36360 26744 36364 26800
rect 36300 26740 36364 26744
rect 36719 26796 36783 26800
rect 36719 26740 36723 26796
rect 36723 26740 36779 26796
rect 36779 26740 36783 26796
rect 36719 26736 36783 26740
rect 36799 26796 36863 26800
rect 36799 26740 36803 26796
rect 36803 26740 36859 26796
rect 36859 26740 36863 26796
rect 36799 26736 36863 26740
rect 36879 26796 36943 26800
rect 36879 26740 36883 26796
rect 36883 26740 36939 26796
rect 36939 26740 36943 26796
rect 36879 26736 36943 26740
rect 36959 26796 37023 26800
rect 36959 26740 36963 26796
rect 36963 26740 37019 26796
rect 37019 26740 37023 26796
rect 36959 26736 37023 26740
rect 37382 26796 37446 26800
rect 37382 26740 37386 26796
rect 37386 26740 37442 26796
rect 37442 26740 37446 26796
rect 37382 26736 37446 26740
rect 37462 26796 37526 26800
rect 37462 26740 37466 26796
rect 37466 26740 37522 26796
rect 37522 26740 37526 26796
rect 37462 26736 37526 26740
rect 37542 26796 37606 26800
rect 37542 26740 37546 26796
rect 37546 26740 37602 26796
rect 37602 26740 37606 26796
rect 37542 26736 37606 26740
rect 37622 26796 37686 26800
rect 37622 26740 37626 26796
rect 37626 26740 37682 26796
rect 37682 26740 37686 26796
rect 37622 26736 37686 26740
rect 35394 26688 35458 26692
rect 35394 26632 35398 26688
rect 35398 26632 35454 26688
rect 35454 26632 35458 26688
rect 35394 26628 35458 26632
rect 35474 26688 35538 26692
rect 35474 26632 35478 26688
rect 35478 26632 35534 26688
rect 35534 26632 35538 26688
rect 35474 26628 35538 26632
rect 35554 26688 35618 26692
rect 35554 26632 35558 26688
rect 35558 26632 35614 26688
rect 35614 26632 35618 26688
rect 35554 26628 35618 26632
rect 35634 26688 35698 26692
rect 35634 26632 35638 26688
rect 35638 26632 35694 26688
rect 35694 26632 35698 26688
rect 35634 26628 35698 26632
rect 36060 26688 36124 26692
rect 36060 26632 36064 26688
rect 36064 26632 36120 26688
rect 36120 26632 36124 26688
rect 36060 26628 36124 26632
rect 36140 26688 36204 26692
rect 36140 26632 36144 26688
rect 36144 26632 36200 26688
rect 36200 26632 36204 26688
rect 36140 26628 36204 26632
rect 36220 26688 36284 26692
rect 36220 26632 36224 26688
rect 36224 26632 36280 26688
rect 36280 26632 36284 26688
rect 36220 26628 36284 26632
rect 36300 26688 36364 26692
rect 36300 26632 36304 26688
rect 36304 26632 36360 26688
rect 36360 26632 36364 26688
rect 36300 26628 36364 26632
rect 36719 26684 36783 26688
rect 36719 26628 36723 26684
rect 36723 26628 36779 26684
rect 36779 26628 36783 26684
rect 36719 26624 36783 26628
rect 36799 26684 36863 26688
rect 36799 26628 36803 26684
rect 36803 26628 36859 26684
rect 36859 26628 36863 26684
rect 36799 26624 36863 26628
rect 36879 26684 36943 26688
rect 36879 26628 36883 26684
rect 36883 26628 36939 26684
rect 36939 26628 36943 26684
rect 36879 26624 36943 26628
rect 36959 26684 37023 26688
rect 36959 26628 36963 26684
rect 36963 26628 37019 26684
rect 37019 26628 37023 26684
rect 36959 26624 37023 26628
rect 37382 26684 37446 26688
rect 37382 26628 37386 26684
rect 37386 26628 37442 26684
rect 37442 26628 37446 26684
rect 37382 26624 37446 26628
rect 37462 26684 37526 26688
rect 37462 26628 37466 26684
rect 37466 26628 37522 26684
rect 37522 26628 37526 26684
rect 37462 26624 37526 26628
rect 37542 26684 37606 26688
rect 37542 26628 37546 26684
rect 37546 26628 37602 26684
rect 37602 26628 37606 26684
rect 37542 26624 37606 26628
rect 37622 26684 37686 26688
rect 37622 26628 37626 26684
rect 37626 26628 37682 26684
rect 37682 26628 37686 26684
rect 37622 26624 37686 26628
rect 35394 26569 35458 26573
rect 35394 26513 35398 26569
rect 35398 26513 35454 26569
rect 35454 26513 35458 26569
rect 35394 26509 35458 26513
rect 35474 26569 35538 26573
rect 35474 26513 35478 26569
rect 35478 26513 35534 26569
rect 35534 26513 35538 26569
rect 35474 26509 35538 26513
rect 35554 26569 35618 26573
rect 35554 26513 35558 26569
rect 35558 26513 35614 26569
rect 35614 26513 35618 26569
rect 35554 26509 35618 26513
rect 35634 26569 35698 26573
rect 35634 26513 35638 26569
rect 35638 26513 35694 26569
rect 35694 26513 35698 26569
rect 35634 26509 35698 26513
rect 36060 26569 36124 26573
rect 36060 26513 36064 26569
rect 36064 26513 36120 26569
rect 36120 26513 36124 26569
rect 36060 26509 36124 26513
rect 36140 26569 36204 26573
rect 36140 26513 36144 26569
rect 36144 26513 36200 26569
rect 36200 26513 36204 26569
rect 36140 26509 36204 26513
rect 36220 26569 36284 26573
rect 36220 26513 36224 26569
rect 36224 26513 36280 26569
rect 36280 26513 36284 26569
rect 36220 26509 36284 26513
rect 36300 26569 36364 26573
rect 36300 26513 36304 26569
rect 36304 26513 36360 26569
rect 36360 26513 36364 26569
rect 36300 26509 36364 26513
rect 36719 26565 36783 26569
rect 36719 26509 36723 26565
rect 36723 26509 36779 26565
rect 36779 26509 36783 26565
rect 36719 26505 36783 26509
rect 36799 26565 36863 26569
rect 36799 26509 36803 26565
rect 36803 26509 36859 26565
rect 36859 26509 36863 26565
rect 36799 26505 36863 26509
rect 36879 26565 36943 26569
rect 36879 26509 36883 26565
rect 36883 26509 36939 26565
rect 36939 26509 36943 26565
rect 36879 26505 36943 26509
rect 36959 26565 37023 26569
rect 36959 26509 36963 26565
rect 36963 26509 37019 26565
rect 37019 26509 37023 26565
rect 36959 26505 37023 26509
rect 37382 26565 37446 26569
rect 37382 26509 37386 26565
rect 37386 26509 37442 26565
rect 37442 26509 37446 26565
rect 37382 26505 37446 26509
rect 37462 26565 37526 26569
rect 37462 26509 37466 26565
rect 37466 26509 37522 26565
rect 37522 26509 37526 26565
rect 37462 26505 37526 26509
rect 37542 26565 37606 26569
rect 37542 26509 37546 26565
rect 37546 26509 37602 26565
rect 37602 26509 37606 26565
rect 37542 26505 37606 26509
rect 37622 26565 37686 26569
rect 37622 26509 37626 26565
rect 37626 26509 37682 26565
rect 37682 26509 37686 26565
rect 37622 26505 37686 26509
rect 46702 26800 46766 26804
rect 46702 26744 46706 26800
rect 46706 26744 46762 26800
rect 46762 26744 46766 26800
rect 46702 26740 46766 26744
rect 46782 26800 46846 26804
rect 46782 26744 46786 26800
rect 46786 26744 46842 26800
rect 46842 26744 46846 26800
rect 46782 26740 46846 26744
rect 46862 26800 46926 26804
rect 46862 26744 46866 26800
rect 46866 26744 46922 26800
rect 46922 26744 46926 26800
rect 46862 26740 46926 26744
rect 46942 26800 47006 26804
rect 46942 26744 46946 26800
rect 46946 26744 47002 26800
rect 47002 26744 47006 26800
rect 46942 26740 47006 26744
rect 47368 26800 47432 26804
rect 47368 26744 47372 26800
rect 47372 26744 47428 26800
rect 47428 26744 47432 26800
rect 47368 26740 47432 26744
rect 47448 26800 47512 26804
rect 47448 26744 47452 26800
rect 47452 26744 47508 26800
rect 47508 26744 47512 26800
rect 47448 26740 47512 26744
rect 47528 26800 47592 26804
rect 47528 26744 47532 26800
rect 47532 26744 47588 26800
rect 47588 26744 47592 26800
rect 47528 26740 47592 26744
rect 47608 26800 47672 26804
rect 47608 26744 47612 26800
rect 47612 26744 47668 26800
rect 47668 26744 47672 26800
rect 47608 26740 47672 26744
rect 48027 26796 48091 26800
rect 48027 26740 48031 26796
rect 48031 26740 48087 26796
rect 48087 26740 48091 26796
rect 48027 26736 48091 26740
rect 48107 26796 48171 26800
rect 48107 26740 48111 26796
rect 48111 26740 48167 26796
rect 48167 26740 48171 26796
rect 48107 26736 48171 26740
rect 48187 26796 48251 26800
rect 48187 26740 48191 26796
rect 48191 26740 48247 26796
rect 48247 26740 48251 26796
rect 48187 26736 48251 26740
rect 48267 26796 48331 26800
rect 48267 26740 48271 26796
rect 48271 26740 48327 26796
rect 48327 26740 48331 26796
rect 48267 26736 48331 26740
rect 48690 26796 48754 26800
rect 48690 26740 48694 26796
rect 48694 26740 48750 26796
rect 48750 26740 48754 26796
rect 48690 26736 48754 26740
rect 48770 26796 48834 26800
rect 48770 26740 48774 26796
rect 48774 26740 48830 26796
rect 48830 26740 48834 26796
rect 48770 26736 48834 26740
rect 48850 26796 48914 26800
rect 48850 26740 48854 26796
rect 48854 26740 48910 26796
rect 48910 26740 48914 26796
rect 48850 26736 48914 26740
rect 48930 26796 48994 26800
rect 48930 26740 48934 26796
rect 48934 26740 48990 26796
rect 48990 26740 48994 26796
rect 48930 26736 48994 26740
rect 46702 26688 46766 26692
rect 46702 26632 46706 26688
rect 46706 26632 46762 26688
rect 46762 26632 46766 26688
rect 46702 26628 46766 26632
rect 46782 26688 46846 26692
rect 46782 26632 46786 26688
rect 46786 26632 46842 26688
rect 46842 26632 46846 26688
rect 46782 26628 46846 26632
rect 46862 26688 46926 26692
rect 46862 26632 46866 26688
rect 46866 26632 46922 26688
rect 46922 26632 46926 26688
rect 46862 26628 46926 26632
rect 46942 26688 47006 26692
rect 46942 26632 46946 26688
rect 46946 26632 47002 26688
rect 47002 26632 47006 26688
rect 46942 26628 47006 26632
rect 47368 26688 47432 26692
rect 47368 26632 47372 26688
rect 47372 26632 47428 26688
rect 47428 26632 47432 26688
rect 47368 26628 47432 26632
rect 47448 26688 47512 26692
rect 47448 26632 47452 26688
rect 47452 26632 47508 26688
rect 47508 26632 47512 26688
rect 47448 26628 47512 26632
rect 47528 26688 47592 26692
rect 47528 26632 47532 26688
rect 47532 26632 47588 26688
rect 47588 26632 47592 26688
rect 47528 26628 47592 26632
rect 47608 26688 47672 26692
rect 47608 26632 47612 26688
rect 47612 26632 47668 26688
rect 47668 26632 47672 26688
rect 47608 26628 47672 26632
rect 48027 26684 48091 26688
rect 48027 26628 48031 26684
rect 48031 26628 48087 26684
rect 48087 26628 48091 26684
rect 48027 26624 48091 26628
rect 48107 26684 48171 26688
rect 48107 26628 48111 26684
rect 48111 26628 48167 26684
rect 48167 26628 48171 26684
rect 48107 26624 48171 26628
rect 48187 26684 48251 26688
rect 48187 26628 48191 26684
rect 48191 26628 48247 26684
rect 48247 26628 48251 26684
rect 48187 26624 48251 26628
rect 48267 26684 48331 26688
rect 48267 26628 48271 26684
rect 48271 26628 48327 26684
rect 48327 26628 48331 26684
rect 48267 26624 48331 26628
rect 48690 26684 48754 26688
rect 48690 26628 48694 26684
rect 48694 26628 48750 26684
rect 48750 26628 48754 26684
rect 48690 26624 48754 26628
rect 48770 26684 48834 26688
rect 48770 26628 48774 26684
rect 48774 26628 48830 26684
rect 48830 26628 48834 26684
rect 48770 26624 48834 26628
rect 48850 26684 48914 26688
rect 48850 26628 48854 26684
rect 48854 26628 48910 26684
rect 48910 26628 48914 26684
rect 48850 26624 48914 26628
rect 48930 26684 48994 26688
rect 48930 26628 48934 26684
rect 48934 26628 48990 26684
rect 48990 26628 48994 26684
rect 48930 26624 48994 26628
rect 46702 26569 46766 26573
rect 46702 26513 46706 26569
rect 46706 26513 46762 26569
rect 46762 26513 46766 26569
rect 46702 26509 46766 26513
rect 46782 26569 46846 26573
rect 46782 26513 46786 26569
rect 46786 26513 46842 26569
rect 46842 26513 46846 26569
rect 46782 26509 46846 26513
rect 46862 26569 46926 26573
rect 46862 26513 46866 26569
rect 46866 26513 46922 26569
rect 46922 26513 46926 26569
rect 46862 26509 46926 26513
rect 46942 26569 47006 26573
rect 46942 26513 46946 26569
rect 46946 26513 47002 26569
rect 47002 26513 47006 26569
rect 46942 26509 47006 26513
rect 47368 26569 47432 26573
rect 47368 26513 47372 26569
rect 47372 26513 47428 26569
rect 47428 26513 47432 26569
rect 47368 26509 47432 26513
rect 47448 26569 47512 26573
rect 47448 26513 47452 26569
rect 47452 26513 47508 26569
rect 47508 26513 47512 26569
rect 47448 26509 47512 26513
rect 47528 26569 47592 26573
rect 47528 26513 47532 26569
rect 47532 26513 47588 26569
rect 47588 26513 47592 26569
rect 47528 26509 47592 26513
rect 47608 26569 47672 26573
rect 47608 26513 47612 26569
rect 47612 26513 47668 26569
rect 47668 26513 47672 26569
rect 47608 26509 47672 26513
rect 48027 26565 48091 26569
rect 48027 26509 48031 26565
rect 48031 26509 48087 26565
rect 48087 26509 48091 26565
rect 48027 26505 48091 26509
rect 48107 26565 48171 26569
rect 48107 26509 48111 26565
rect 48111 26509 48167 26565
rect 48167 26509 48171 26565
rect 48107 26505 48171 26509
rect 48187 26565 48251 26569
rect 48187 26509 48191 26565
rect 48191 26509 48247 26565
rect 48247 26509 48251 26565
rect 48187 26505 48251 26509
rect 48267 26565 48331 26569
rect 48267 26509 48271 26565
rect 48271 26509 48327 26565
rect 48327 26509 48331 26565
rect 48267 26505 48331 26509
rect 48690 26565 48754 26569
rect 48690 26509 48694 26565
rect 48694 26509 48750 26565
rect 48750 26509 48754 26565
rect 48690 26505 48754 26509
rect 48770 26565 48834 26569
rect 48770 26509 48774 26565
rect 48774 26509 48830 26565
rect 48830 26509 48834 26565
rect 48770 26505 48834 26509
rect 48850 26565 48914 26569
rect 48850 26509 48854 26565
rect 48854 26509 48910 26565
rect 48910 26509 48914 26565
rect 48850 26505 48914 26509
rect 48930 26565 48994 26569
rect 48930 26509 48934 26565
rect 48934 26509 48990 26565
rect 48990 26509 48994 26565
rect 48930 26505 48994 26509
rect 50831 26800 50895 26804
rect 50831 26744 50835 26800
rect 50835 26744 50891 26800
rect 50891 26744 50895 26800
rect 50831 26740 50895 26744
rect 50911 26800 50975 26804
rect 50911 26744 50915 26800
rect 50915 26744 50971 26800
rect 50971 26744 50975 26800
rect 50911 26740 50975 26744
rect 50991 26800 51055 26804
rect 50991 26744 50995 26800
rect 50995 26744 51051 26800
rect 51051 26744 51055 26800
rect 50991 26740 51055 26744
rect 51071 26800 51135 26804
rect 51071 26744 51075 26800
rect 51075 26744 51131 26800
rect 51131 26744 51135 26800
rect 51071 26740 51135 26744
rect 51497 26800 51561 26804
rect 51497 26744 51501 26800
rect 51501 26744 51557 26800
rect 51557 26744 51561 26800
rect 51497 26740 51561 26744
rect 51577 26800 51641 26804
rect 51577 26744 51581 26800
rect 51581 26744 51637 26800
rect 51637 26744 51641 26800
rect 51577 26740 51641 26744
rect 51657 26800 51721 26804
rect 51657 26744 51661 26800
rect 51661 26744 51717 26800
rect 51717 26744 51721 26800
rect 51657 26740 51721 26744
rect 51737 26800 51801 26804
rect 51737 26744 51741 26800
rect 51741 26744 51797 26800
rect 51797 26744 51801 26800
rect 51737 26740 51801 26744
rect 52156 26796 52220 26800
rect 52156 26740 52160 26796
rect 52160 26740 52216 26796
rect 52216 26740 52220 26796
rect 52156 26736 52220 26740
rect 52236 26796 52300 26800
rect 52236 26740 52240 26796
rect 52240 26740 52296 26796
rect 52296 26740 52300 26796
rect 52236 26736 52300 26740
rect 52316 26796 52380 26800
rect 52316 26740 52320 26796
rect 52320 26740 52376 26796
rect 52376 26740 52380 26796
rect 52316 26736 52380 26740
rect 52396 26796 52460 26800
rect 52396 26740 52400 26796
rect 52400 26740 52456 26796
rect 52456 26740 52460 26796
rect 52396 26736 52460 26740
rect 52819 26796 52883 26800
rect 52819 26740 52823 26796
rect 52823 26740 52879 26796
rect 52879 26740 52883 26796
rect 52819 26736 52883 26740
rect 52899 26796 52963 26800
rect 52899 26740 52903 26796
rect 52903 26740 52959 26796
rect 52959 26740 52963 26796
rect 52899 26736 52963 26740
rect 52979 26796 53043 26800
rect 52979 26740 52983 26796
rect 52983 26740 53039 26796
rect 53039 26740 53043 26796
rect 52979 26736 53043 26740
rect 53059 26796 53123 26800
rect 53059 26740 53063 26796
rect 53063 26740 53119 26796
rect 53119 26740 53123 26796
rect 53059 26736 53123 26740
rect 50831 26688 50895 26692
rect 50831 26632 50835 26688
rect 50835 26632 50891 26688
rect 50891 26632 50895 26688
rect 50831 26628 50895 26632
rect 50911 26688 50975 26692
rect 50911 26632 50915 26688
rect 50915 26632 50971 26688
rect 50971 26632 50975 26688
rect 50911 26628 50975 26632
rect 50991 26688 51055 26692
rect 50991 26632 50995 26688
rect 50995 26632 51051 26688
rect 51051 26632 51055 26688
rect 50991 26628 51055 26632
rect 51071 26688 51135 26692
rect 51071 26632 51075 26688
rect 51075 26632 51131 26688
rect 51131 26632 51135 26688
rect 51071 26628 51135 26632
rect 51497 26688 51561 26692
rect 51497 26632 51501 26688
rect 51501 26632 51557 26688
rect 51557 26632 51561 26688
rect 51497 26628 51561 26632
rect 51577 26688 51641 26692
rect 51577 26632 51581 26688
rect 51581 26632 51637 26688
rect 51637 26632 51641 26688
rect 51577 26628 51641 26632
rect 51657 26688 51721 26692
rect 51657 26632 51661 26688
rect 51661 26632 51717 26688
rect 51717 26632 51721 26688
rect 51657 26628 51721 26632
rect 51737 26688 51801 26692
rect 51737 26632 51741 26688
rect 51741 26632 51797 26688
rect 51797 26632 51801 26688
rect 51737 26628 51801 26632
rect 52156 26684 52220 26688
rect 52156 26628 52160 26684
rect 52160 26628 52216 26684
rect 52216 26628 52220 26684
rect 52156 26624 52220 26628
rect 52236 26684 52300 26688
rect 52236 26628 52240 26684
rect 52240 26628 52296 26684
rect 52296 26628 52300 26684
rect 52236 26624 52300 26628
rect 52316 26684 52380 26688
rect 52316 26628 52320 26684
rect 52320 26628 52376 26684
rect 52376 26628 52380 26684
rect 52316 26624 52380 26628
rect 52396 26684 52460 26688
rect 52396 26628 52400 26684
rect 52400 26628 52456 26684
rect 52456 26628 52460 26684
rect 52396 26624 52460 26628
rect 52819 26684 52883 26688
rect 52819 26628 52823 26684
rect 52823 26628 52879 26684
rect 52879 26628 52883 26684
rect 52819 26624 52883 26628
rect 52899 26684 52963 26688
rect 52899 26628 52903 26684
rect 52903 26628 52959 26684
rect 52959 26628 52963 26684
rect 52899 26624 52963 26628
rect 52979 26684 53043 26688
rect 52979 26628 52983 26684
rect 52983 26628 53039 26684
rect 53039 26628 53043 26684
rect 52979 26624 53043 26628
rect 53059 26684 53123 26688
rect 53059 26628 53063 26684
rect 53063 26628 53119 26684
rect 53119 26628 53123 26684
rect 53059 26624 53123 26628
rect 50831 26569 50895 26573
rect 50831 26513 50835 26569
rect 50835 26513 50891 26569
rect 50891 26513 50895 26569
rect 50831 26509 50895 26513
rect 50911 26569 50975 26573
rect 50911 26513 50915 26569
rect 50915 26513 50971 26569
rect 50971 26513 50975 26569
rect 50911 26509 50975 26513
rect 50991 26569 51055 26573
rect 50991 26513 50995 26569
rect 50995 26513 51051 26569
rect 51051 26513 51055 26569
rect 50991 26509 51055 26513
rect 51071 26569 51135 26573
rect 51071 26513 51075 26569
rect 51075 26513 51131 26569
rect 51131 26513 51135 26569
rect 51071 26509 51135 26513
rect 51497 26569 51561 26573
rect 51497 26513 51501 26569
rect 51501 26513 51557 26569
rect 51557 26513 51561 26569
rect 51497 26509 51561 26513
rect 51577 26569 51641 26573
rect 51577 26513 51581 26569
rect 51581 26513 51637 26569
rect 51637 26513 51641 26569
rect 51577 26509 51641 26513
rect 51657 26569 51721 26573
rect 51657 26513 51661 26569
rect 51661 26513 51717 26569
rect 51717 26513 51721 26569
rect 51657 26509 51721 26513
rect 51737 26569 51801 26573
rect 51737 26513 51741 26569
rect 51741 26513 51797 26569
rect 51797 26513 51801 26569
rect 51737 26509 51801 26513
rect 52156 26565 52220 26569
rect 52156 26509 52160 26565
rect 52160 26509 52216 26565
rect 52216 26509 52220 26565
rect 52156 26505 52220 26509
rect 52236 26565 52300 26569
rect 52236 26509 52240 26565
rect 52240 26509 52296 26565
rect 52296 26509 52300 26565
rect 52236 26505 52300 26509
rect 52316 26565 52380 26569
rect 52316 26509 52320 26565
rect 52320 26509 52376 26565
rect 52376 26509 52380 26565
rect 52316 26505 52380 26509
rect 52396 26565 52460 26569
rect 52396 26509 52400 26565
rect 52400 26509 52456 26565
rect 52456 26509 52460 26565
rect 52396 26505 52460 26509
rect 52819 26565 52883 26569
rect 52819 26509 52823 26565
rect 52823 26509 52879 26565
rect 52879 26509 52883 26565
rect 52819 26505 52883 26509
rect 52899 26565 52963 26569
rect 52899 26509 52903 26565
rect 52903 26509 52959 26565
rect 52959 26509 52963 26565
rect 52899 26505 52963 26509
rect 52979 26565 53043 26569
rect 52979 26509 52983 26565
rect 52983 26509 53039 26565
rect 53039 26509 53043 26565
rect 52979 26505 53043 26509
rect 53059 26565 53123 26569
rect 53059 26509 53063 26565
rect 53063 26509 53119 26565
rect 53119 26509 53123 26565
rect 53059 26505 53123 26509
rect 40315 13620 40379 13624
rect 40315 13564 40319 13620
rect 40319 13564 40375 13620
rect 40375 13564 40379 13620
rect 40315 13560 40379 13564
rect 40395 13620 40459 13624
rect 40395 13564 40399 13620
rect 40399 13564 40455 13620
rect 40455 13564 40459 13620
rect 40395 13560 40459 13564
rect 40315 13501 40379 13505
rect 40315 13445 40319 13501
rect 40319 13445 40375 13501
rect 40375 13445 40379 13501
rect 40315 13441 40379 13445
rect 40395 13501 40459 13505
rect 40395 13445 40399 13501
rect 40399 13445 40455 13501
rect 40455 13445 40459 13501
rect 40395 13441 40459 13445
rect 40315 13380 40379 13384
rect 40315 13324 40319 13380
rect 40319 13324 40375 13380
rect 40375 13324 40379 13380
rect 40315 13320 40379 13324
rect 40395 13380 40459 13384
rect 40395 13324 40399 13380
rect 40399 13324 40455 13380
rect 40455 13324 40459 13380
rect 40395 13320 40459 13324
rect 40315 13273 40379 13277
rect 40315 13217 40319 13273
rect 40319 13217 40375 13273
rect 40375 13217 40379 13273
rect 40315 13213 40379 13217
rect 40395 13273 40459 13277
rect 40395 13217 40399 13273
rect 40399 13217 40455 13273
rect 40455 13217 40459 13273
rect 40395 13213 40459 13217
rect 31265 13108 31329 13112
rect 31265 13052 31269 13108
rect 31269 13052 31325 13108
rect 31325 13052 31329 13108
rect 31265 13048 31329 13052
rect 31345 13108 31409 13112
rect 31345 13052 31349 13108
rect 31349 13052 31405 13108
rect 31405 13052 31409 13108
rect 31345 13048 31409 13052
rect 31425 13108 31489 13112
rect 31425 13052 31429 13108
rect 31429 13052 31485 13108
rect 31485 13052 31489 13108
rect 31425 13048 31489 13052
rect 31505 13108 31569 13112
rect 31505 13052 31509 13108
rect 31509 13052 31565 13108
rect 31565 13052 31569 13108
rect 31505 13048 31569 13052
rect 31931 13108 31995 13112
rect 31931 13052 31935 13108
rect 31935 13052 31991 13108
rect 31991 13052 31995 13108
rect 31931 13048 31995 13052
rect 32011 13108 32075 13112
rect 32011 13052 32015 13108
rect 32015 13052 32071 13108
rect 32071 13052 32075 13108
rect 32011 13048 32075 13052
rect 32091 13108 32155 13112
rect 32091 13052 32095 13108
rect 32095 13052 32151 13108
rect 32151 13052 32155 13108
rect 32091 13048 32155 13052
rect 32171 13108 32235 13112
rect 32171 13052 32175 13108
rect 32175 13052 32231 13108
rect 32231 13052 32235 13108
rect 32171 13048 32235 13052
rect 32590 13104 32654 13108
rect 32590 13048 32594 13104
rect 32594 13048 32650 13104
rect 32650 13048 32654 13104
rect 32590 13044 32654 13048
rect 32670 13104 32734 13108
rect 32670 13048 32674 13104
rect 32674 13048 32730 13104
rect 32730 13048 32734 13104
rect 32670 13044 32734 13048
rect 32750 13104 32814 13108
rect 32750 13048 32754 13104
rect 32754 13048 32810 13104
rect 32810 13048 32814 13104
rect 32750 13044 32814 13048
rect 32830 13104 32894 13108
rect 32830 13048 32834 13104
rect 32834 13048 32890 13104
rect 32890 13048 32894 13104
rect 32830 13044 32894 13048
rect 33253 13104 33317 13108
rect 33253 13048 33257 13104
rect 33257 13048 33313 13104
rect 33313 13048 33317 13104
rect 33253 13044 33317 13048
rect 33333 13104 33397 13108
rect 33333 13048 33337 13104
rect 33337 13048 33393 13104
rect 33393 13048 33397 13104
rect 33333 13044 33397 13048
rect 33413 13104 33477 13108
rect 33413 13048 33417 13104
rect 33417 13048 33473 13104
rect 33473 13048 33477 13104
rect 33413 13044 33477 13048
rect 33493 13104 33557 13108
rect 33493 13048 33497 13104
rect 33497 13048 33553 13104
rect 33553 13048 33557 13104
rect 33493 13044 33557 13048
rect 31265 12996 31329 13000
rect 31265 12940 31269 12996
rect 31269 12940 31325 12996
rect 31325 12940 31329 12996
rect 31265 12936 31329 12940
rect 31345 12996 31409 13000
rect 31345 12940 31349 12996
rect 31349 12940 31405 12996
rect 31405 12940 31409 12996
rect 31345 12936 31409 12940
rect 31425 12996 31489 13000
rect 31425 12940 31429 12996
rect 31429 12940 31485 12996
rect 31485 12940 31489 12996
rect 31425 12936 31489 12940
rect 31505 12996 31569 13000
rect 31505 12940 31509 12996
rect 31509 12940 31565 12996
rect 31565 12940 31569 12996
rect 31505 12936 31569 12940
rect 31931 12996 31995 13000
rect 31931 12940 31935 12996
rect 31935 12940 31991 12996
rect 31991 12940 31995 12996
rect 31931 12936 31995 12940
rect 32011 12996 32075 13000
rect 32011 12940 32015 12996
rect 32015 12940 32071 12996
rect 32071 12940 32075 12996
rect 32011 12936 32075 12940
rect 32091 12996 32155 13000
rect 32091 12940 32095 12996
rect 32095 12940 32151 12996
rect 32151 12940 32155 12996
rect 32091 12936 32155 12940
rect 32171 12996 32235 13000
rect 32171 12940 32175 12996
rect 32175 12940 32231 12996
rect 32231 12940 32235 12996
rect 32171 12936 32235 12940
rect 32590 12992 32654 12996
rect 32590 12936 32594 12992
rect 32594 12936 32650 12992
rect 32650 12936 32654 12992
rect 32590 12932 32654 12936
rect 32670 12992 32734 12996
rect 32670 12936 32674 12992
rect 32674 12936 32730 12992
rect 32730 12936 32734 12992
rect 32670 12932 32734 12936
rect 32750 12992 32814 12996
rect 32750 12936 32754 12992
rect 32754 12936 32810 12992
rect 32810 12936 32814 12992
rect 32750 12932 32814 12936
rect 32830 12992 32894 12996
rect 32830 12936 32834 12992
rect 32834 12936 32890 12992
rect 32890 12936 32894 12992
rect 32830 12932 32894 12936
rect 33253 12992 33317 12996
rect 33253 12936 33257 12992
rect 33257 12936 33313 12992
rect 33313 12936 33317 12992
rect 33253 12932 33317 12936
rect 33333 12992 33397 12996
rect 33333 12936 33337 12992
rect 33337 12936 33393 12992
rect 33393 12936 33397 12992
rect 33333 12932 33397 12936
rect 33413 12992 33477 12996
rect 33413 12936 33417 12992
rect 33417 12936 33473 12992
rect 33473 12936 33477 12992
rect 33413 12932 33477 12936
rect 33493 12992 33557 12996
rect 33493 12936 33497 12992
rect 33497 12936 33553 12992
rect 33553 12936 33557 12992
rect 33493 12932 33557 12936
rect 31265 12877 31329 12881
rect 31265 12821 31269 12877
rect 31269 12821 31325 12877
rect 31325 12821 31329 12877
rect 31265 12817 31329 12821
rect 31345 12877 31409 12881
rect 31345 12821 31349 12877
rect 31349 12821 31405 12877
rect 31405 12821 31409 12877
rect 31345 12817 31409 12821
rect 31425 12877 31489 12881
rect 31425 12821 31429 12877
rect 31429 12821 31485 12877
rect 31485 12821 31489 12877
rect 31425 12817 31489 12821
rect 31505 12877 31569 12881
rect 31505 12821 31509 12877
rect 31509 12821 31565 12877
rect 31565 12821 31569 12877
rect 31505 12817 31569 12821
rect 31931 12877 31995 12881
rect 31931 12821 31935 12877
rect 31935 12821 31991 12877
rect 31991 12821 31995 12877
rect 31931 12817 31995 12821
rect 32011 12877 32075 12881
rect 32011 12821 32015 12877
rect 32015 12821 32071 12877
rect 32071 12821 32075 12877
rect 32011 12817 32075 12821
rect 32091 12877 32155 12881
rect 32091 12821 32095 12877
rect 32095 12821 32151 12877
rect 32151 12821 32155 12877
rect 32091 12817 32155 12821
rect 32171 12877 32235 12881
rect 32171 12821 32175 12877
rect 32175 12821 32231 12877
rect 32231 12821 32235 12877
rect 32171 12817 32235 12821
rect 32590 12873 32654 12877
rect 32590 12817 32594 12873
rect 32594 12817 32650 12873
rect 32650 12817 32654 12873
rect 32590 12813 32654 12817
rect 32670 12873 32734 12877
rect 32670 12817 32674 12873
rect 32674 12817 32730 12873
rect 32730 12817 32734 12873
rect 32670 12813 32734 12817
rect 32750 12873 32814 12877
rect 32750 12817 32754 12873
rect 32754 12817 32810 12873
rect 32810 12817 32814 12873
rect 32750 12813 32814 12817
rect 32830 12873 32894 12877
rect 32830 12817 32834 12873
rect 32834 12817 32890 12873
rect 32890 12817 32894 12873
rect 32830 12813 32894 12817
rect 33253 12873 33317 12877
rect 33253 12817 33257 12873
rect 33257 12817 33313 12873
rect 33313 12817 33317 12873
rect 33253 12813 33317 12817
rect 33333 12873 33397 12877
rect 33333 12817 33337 12873
rect 33337 12817 33393 12873
rect 33393 12817 33397 12873
rect 33333 12813 33397 12817
rect 33413 12873 33477 12877
rect 33413 12817 33417 12873
rect 33417 12817 33473 12873
rect 33473 12817 33477 12873
rect 33413 12813 33477 12817
rect 33493 12873 33557 12877
rect 33493 12817 33497 12873
rect 33497 12817 33553 12873
rect 33553 12817 33557 12873
rect 33493 12813 33557 12817
rect 35394 13108 35458 13112
rect 35394 13052 35398 13108
rect 35398 13052 35454 13108
rect 35454 13052 35458 13108
rect 35394 13048 35458 13052
rect 35474 13108 35538 13112
rect 35474 13052 35478 13108
rect 35478 13052 35534 13108
rect 35534 13052 35538 13108
rect 35474 13048 35538 13052
rect 35554 13108 35618 13112
rect 35554 13052 35558 13108
rect 35558 13052 35614 13108
rect 35614 13052 35618 13108
rect 35554 13048 35618 13052
rect 35634 13108 35698 13112
rect 35634 13052 35638 13108
rect 35638 13052 35694 13108
rect 35694 13052 35698 13108
rect 35634 13048 35698 13052
rect 36060 13108 36124 13112
rect 36060 13052 36064 13108
rect 36064 13052 36120 13108
rect 36120 13052 36124 13108
rect 36060 13048 36124 13052
rect 36140 13108 36204 13112
rect 36140 13052 36144 13108
rect 36144 13052 36200 13108
rect 36200 13052 36204 13108
rect 36140 13048 36204 13052
rect 36220 13108 36284 13112
rect 36220 13052 36224 13108
rect 36224 13052 36280 13108
rect 36280 13052 36284 13108
rect 36220 13048 36284 13052
rect 36300 13108 36364 13112
rect 36300 13052 36304 13108
rect 36304 13052 36360 13108
rect 36360 13052 36364 13108
rect 36300 13048 36364 13052
rect 36719 13104 36783 13108
rect 36719 13048 36723 13104
rect 36723 13048 36779 13104
rect 36779 13048 36783 13104
rect 36719 13044 36783 13048
rect 36799 13104 36863 13108
rect 36799 13048 36803 13104
rect 36803 13048 36859 13104
rect 36859 13048 36863 13104
rect 36799 13044 36863 13048
rect 36879 13104 36943 13108
rect 36879 13048 36883 13104
rect 36883 13048 36939 13104
rect 36939 13048 36943 13104
rect 36879 13044 36943 13048
rect 36959 13104 37023 13108
rect 36959 13048 36963 13104
rect 36963 13048 37019 13104
rect 37019 13048 37023 13104
rect 36959 13044 37023 13048
rect 37382 13104 37446 13108
rect 37382 13048 37386 13104
rect 37386 13048 37442 13104
rect 37442 13048 37446 13104
rect 37382 13044 37446 13048
rect 37462 13104 37526 13108
rect 37462 13048 37466 13104
rect 37466 13048 37522 13104
rect 37522 13048 37526 13104
rect 37462 13044 37526 13048
rect 37542 13104 37606 13108
rect 37542 13048 37546 13104
rect 37546 13048 37602 13104
rect 37602 13048 37606 13104
rect 37542 13044 37606 13048
rect 37622 13104 37686 13108
rect 37622 13048 37626 13104
rect 37626 13048 37682 13104
rect 37682 13048 37686 13104
rect 37622 13044 37686 13048
rect 35394 12996 35458 13000
rect 35394 12940 35398 12996
rect 35398 12940 35454 12996
rect 35454 12940 35458 12996
rect 35394 12936 35458 12940
rect 35474 12996 35538 13000
rect 35474 12940 35478 12996
rect 35478 12940 35534 12996
rect 35534 12940 35538 12996
rect 35474 12936 35538 12940
rect 35554 12996 35618 13000
rect 35554 12940 35558 12996
rect 35558 12940 35614 12996
rect 35614 12940 35618 12996
rect 35554 12936 35618 12940
rect 35634 12996 35698 13000
rect 35634 12940 35638 12996
rect 35638 12940 35694 12996
rect 35694 12940 35698 12996
rect 35634 12936 35698 12940
rect 36060 12996 36124 13000
rect 36060 12940 36064 12996
rect 36064 12940 36120 12996
rect 36120 12940 36124 12996
rect 36060 12936 36124 12940
rect 36140 12996 36204 13000
rect 36140 12940 36144 12996
rect 36144 12940 36200 12996
rect 36200 12940 36204 12996
rect 36140 12936 36204 12940
rect 36220 12996 36284 13000
rect 36220 12940 36224 12996
rect 36224 12940 36280 12996
rect 36280 12940 36284 12996
rect 36220 12936 36284 12940
rect 36300 12996 36364 13000
rect 36300 12940 36304 12996
rect 36304 12940 36360 12996
rect 36360 12940 36364 12996
rect 36300 12936 36364 12940
rect 36719 12992 36783 12996
rect 36719 12936 36723 12992
rect 36723 12936 36779 12992
rect 36779 12936 36783 12992
rect 36719 12932 36783 12936
rect 36799 12992 36863 12996
rect 36799 12936 36803 12992
rect 36803 12936 36859 12992
rect 36859 12936 36863 12992
rect 36799 12932 36863 12936
rect 36879 12992 36943 12996
rect 36879 12936 36883 12992
rect 36883 12936 36939 12992
rect 36939 12936 36943 12992
rect 36879 12932 36943 12936
rect 36959 12992 37023 12996
rect 36959 12936 36963 12992
rect 36963 12936 37019 12992
rect 37019 12936 37023 12992
rect 36959 12932 37023 12936
rect 37382 12992 37446 12996
rect 37382 12936 37386 12992
rect 37386 12936 37442 12992
rect 37442 12936 37446 12992
rect 37382 12932 37446 12936
rect 37462 12992 37526 12996
rect 37462 12936 37466 12992
rect 37466 12936 37522 12992
rect 37522 12936 37526 12992
rect 37462 12932 37526 12936
rect 37542 12992 37606 12996
rect 37542 12936 37546 12992
rect 37546 12936 37602 12992
rect 37602 12936 37606 12992
rect 37542 12932 37606 12936
rect 37622 12992 37686 12996
rect 37622 12936 37626 12992
rect 37626 12936 37682 12992
rect 37682 12936 37686 12992
rect 37622 12932 37686 12936
rect 35394 12877 35458 12881
rect 35394 12821 35398 12877
rect 35398 12821 35454 12877
rect 35454 12821 35458 12877
rect 35394 12817 35458 12821
rect 35474 12877 35538 12881
rect 35474 12821 35478 12877
rect 35478 12821 35534 12877
rect 35534 12821 35538 12877
rect 35474 12817 35538 12821
rect 35554 12877 35618 12881
rect 35554 12821 35558 12877
rect 35558 12821 35614 12877
rect 35614 12821 35618 12877
rect 35554 12817 35618 12821
rect 35634 12877 35698 12881
rect 35634 12821 35638 12877
rect 35638 12821 35694 12877
rect 35694 12821 35698 12877
rect 35634 12817 35698 12821
rect 36060 12877 36124 12881
rect 36060 12821 36064 12877
rect 36064 12821 36120 12877
rect 36120 12821 36124 12877
rect 36060 12817 36124 12821
rect 36140 12877 36204 12881
rect 36140 12821 36144 12877
rect 36144 12821 36200 12877
rect 36200 12821 36204 12877
rect 36140 12817 36204 12821
rect 36220 12877 36284 12881
rect 36220 12821 36224 12877
rect 36224 12821 36280 12877
rect 36280 12821 36284 12877
rect 36220 12817 36284 12821
rect 36300 12877 36364 12881
rect 36300 12821 36304 12877
rect 36304 12821 36360 12877
rect 36360 12821 36364 12877
rect 36300 12817 36364 12821
rect 36719 12873 36783 12877
rect 36719 12817 36723 12873
rect 36723 12817 36779 12873
rect 36779 12817 36783 12873
rect 36719 12813 36783 12817
rect 36799 12873 36863 12877
rect 36799 12817 36803 12873
rect 36803 12817 36859 12873
rect 36859 12817 36863 12873
rect 36799 12813 36863 12817
rect 36879 12873 36943 12877
rect 36879 12817 36883 12873
rect 36883 12817 36939 12873
rect 36939 12817 36943 12873
rect 36879 12813 36943 12817
rect 36959 12873 37023 12877
rect 36959 12817 36963 12873
rect 36963 12817 37019 12873
rect 37019 12817 37023 12873
rect 36959 12813 37023 12817
rect 37382 12873 37446 12877
rect 37382 12817 37386 12873
rect 37386 12817 37442 12873
rect 37442 12817 37446 12873
rect 37382 12813 37446 12817
rect 37462 12873 37526 12877
rect 37462 12817 37466 12873
rect 37466 12817 37522 12873
rect 37522 12817 37526 12873
rect 37462 12813 37526 12817
rect 37542 12873 37606 12877
rect 37542 12817 37546 12873
rect 37546 12817 37602 12873
rect 37602 12817 37606 12873
rect 37542 12813 37606 12817
rect 37622 12873 37686 12877
rect 37622 12817 37626 12873
rect 37626 12817 37682 12873
rect 37682 12817 37686 12873
rect 37622 12813 37686 12817
rect 40315 13147 40379 13151
rect 40315 13091 40319 13147
rect 40319 13091 40375 13147
rect 40375 13091 40379 13147
rect 40315 13087 40379 13091
rect 40395 13147 40459 13151
rect 40395 13091 40399 13147
rect 40399 13091 40455 13147
rect 40455 13091 40459 13147
rect 40395 13087 40459 13091
rect 40315 13035 40379 13039
rect 40315 12979 40319 13035
rect 40319 12979 40375 13035
rect 40375 12979 40379 13035
rect 40315 12975 40379 12979
rect 40395 13035 40459 13039
rect 40395 12979 40399 13035
rect 40399 12979 40455 13035
rect 40455 12979 40459 13035
rect 40395 12975 40459 12979
rect 40315 12916 40379 12920
rect 40315 12860 40319 12916
rect 40319 12860 40375 12916
rect 40375 12860 40379 12916
rect 40315 12856 40379 12860
rect 40395 12916 40459 12920
rect 40395 12860 40399 12916
rect 40399 12860 40455 12916
rect 40455 12860 40459 12916
rect 40395 12856 40459 12860
rect 42790 13564 42854 13568
rect 42790 13508 42794 13564
rect 42794 13508 42850 13564
rect 42850 13508 42854 13564
rect 42790 13504 42854 13508
rect 42870 13564 42934 13568
rect 42870 13508 42874 13564
rect 42874 13508 42930 13564
rect 42930 13508 42934 13564
rect 42870 13504 42934 13508
rect 42790 13441 42854 13445
rect 42790 13385 42794 13441
rect 42794 13385 42850 13441
rect 42850 13385 42854 13441
rect 42790 13381 42854 13385
rect 42870 13441 42934 13445
rect 42870 13385 42874 13441
rect 42874 13385 42930 13441
rect 42930 13385 42934 13441
rect 42870 13381 42934 13385
rect 42790 13329 42854 13333
rect 42790 13273 42794 13329
rect 42794 13273 42850 13329
rect 42850 13273 42854 13329
rect 42790 13269 42854 13273
rect 42870 13329 42934 13333
rect 42870 13273 42874 13329
rect 42874 13273 42930 13329
rect 42930 13273 42934 13329
rect 42870 13269 42934 13273
rect 42790 13210 42854 13214
rect 42790 13154 42794 13210
rect 42794 13154 42850 13210
rect 42850 13154 42854 13210
rect 42790 13150 42854 13154
rect 42870 13210 42934 13214
rect 42870 13154 42874 13210
rect 42874 13154 42930 13210
rect 42930 13154 42934 13210
rect 42870 13150 42934 13154
rect 42790 13086 42854 13090
rect 42790 13030 42794 13086
rect 42794 13030 42850 13086
rect 42850 13030 42854 13086
rect 42790 13026 42854 13030
rect 42870 13086 42934 13090
rect 42870 13030 42874 13086
rect 42874 13030 42930 13086
rect 42930 13030 42934 13086
rect 42870 13026 42934 13030
rect 42790 12979 42854 12983
rect 42790 12923 42794 12979
rect 42794 12923 42850 12979
rect 42850 12923 42854 12979
rect 42790 12919 42854 12923
rect 42870 12979 42934 12983
rect 42870 12923 42874 12979
rect 42874 12923 42930 12979
rect 42930 12923 42934 12979
rect 42870 12919 42934 12923
rect 46702 13108 46766 13112
rect 46702 13052 46706 13108
rect 46706 13052 46762 13108
rect 46762 13052 46766 13108
rect 46702 13048 46766 13052
rect 46782 13108 46846 13112
rect 46782 13052 46786 13108
rect 46786 13052 46842 13108
rect 46842 13052 46846 13108
rect 46782 13048 46846 13052
rect 46862 13108 46926 13112
rect 46862 13052 46866 13108
rect 46866 13052 46922 13108
rect 46922 13052 46926 13108
rect 46862 13048 46926 13052
rect 46942 13108 47006 13112
rect 46942 13052 46946 13108
rect 46946 13052 47002 13108
rect 47002 13052 47006 13108
rect 46942 13048 47006 13052
rect 47368 13108 47432 13112
rect 47368 13052 47372 13108
rect 47372 13052 47428 13108
rect 47428 13052 47432 13108
rect 47368 13048 47432 13052
rect 47448 13108 47512 13112
rect 47448 13052 47452 13108
rect 47452 13052 47508 13108
rect 47508 13052 47512 13108
rect 47448 13048 47512 13052
rect 47528 13108 47592 13112
rect 47528 13052 47532 13108
rect 47532 13052 47588 13108
rect 47588 13052 47592 13108
rect 47528 13048 47592 13052
rect 47608 13108 47672 13112
rect 47608 13052 47612 13108
rect 47612 13052 47668 13108
rect 47668 13052 47672 13108
rect 47608 13048 47672 13052
rect 48027 13104 48091 13108
rect 48027 13048 48031 13104
rect 48031 13048 48087 13104
rect 48087 13048 48091 13104
rect 48027 13044 48091 13048
rect 48107 13104 48171 13108
rect 48107 13048 48111 13104
rect 48111 13048 48167 13104
rect 48167 13048 48171 13104
rect 48107 13044 48171 13048
rect 48187 13104 48251 13108
rect 48187 13048 48191 13104
rect 48191 13048 48247 13104
rect 48247 13048 48251 13104
rect 48187 13044 48251 13048
rect 48267 13104 48331 13108
rect 48267 13048 48271 13104
rect 48271 13048 48327 13104
rect 48327 13048 48331 13104
rect 48267 13044 48331 13048
rect 48690 13104 48754 13108
rect 48690 13048 48694 13104
rect 48694 13048 48750 13104
rect 48750 13048 48754 13104
rect 48690 13044 48754 13048
rect 48770 13104 48834 13108
rect 48770 13048 48774 13104
rect 48774 13048 48830 13104
rect 48830 13048 48834 13104
rect 48770 13044 48834 13048
rect 48850 13104 48914 13108
rect 48850 13048 48854 13104
rect 48854 13048 48910 13104
rect 48910 13048 48914 13104
rect 48850 13044 48914 13048
rect 48930 13104 48994 13108
rect 48930 13048 48934 13104
rect 48934 13048 48990 13104
rect 48990 13048 48994 13104
rect 48930 13044 48994 13048
rect 46702 12996 46766 13000
rect 46702 12940 46706 12996
rect 46706 12940 46762 12996
rect 46762 12940 46766 12996
rect 46702 12936 46766 12940
rect 46782 12996 46846 13000
rect 46782 12940 46786 12996
rect 46786 12940 46842 12996
rect 46842 12940 46846 12996
rect 46782 12936 46846 12940
rect 46862 12996 46926 13000
rect 46862 12940 46866 12996
rect 46866 12940 46922 12996
rect 46922 12940 46926 12996
rect 46862 12936 46926 12940
rect 46942 12996 47006 13000
rect 46942 12940 46946 12996
rect 46946 12940 47002 12996
rect 47002 12940 47006 12996
rect 46942 12936 47006 12940
rect 47368 12996 47432 13000
rect 47368 12940 47372 12996
rect 47372 12940 47428 12996
rect 47428 12940 47432 12996
rect 47368 12936 47432 12940
rect 47448 12996 47512 13000
rect 47448 12940 47452 12996
rect 47452 12940 47508 12996
rect 47508 12940 47512 12996
rect 47448 12936 47512 12940
rect 47528 12996 47592 13000
rect 47528 12940 47532 12996
rect 47532 12940 47588 12996
rect 47588 12940 47592 12996
rect 47528 12936 47592 12940
rect 47608 12996 47672 13000
rect 47608 12940 47612 12996
rect 47612 12940 47668 12996
rect 47668 12940 47672 12996
rect 47608 12936 47672 12940
rect 48027 12992 48091 12996
rect 48027 12936 48031 12992
rect 48031 12936 48087 12992
rect 48087 12936 48091 12992
rect 48027 12932 48091 12936
rect 48107 12992 48171 12996
rect 48107 12936 48111 12992
rect 48111 12936 48167 12992
rect 48167 12936 48171 12992
rect 48107 12932 48171 12936
rect 48187 12992 48251 12996
rect 48187 12936 48191 12992
rect 48191 12936 48247 12992
rect 48247 12936 48251 12992
rect 48187 12932 48251 12936
rect 48267 12992 48331 12996
rect 48267 12936 48271 12992
rect 48271 12936 48327 12992
rect 48327 12936 48331 12992
rect 48267 12932 48331 12936
rect 48690 12992 48754 12996
rect 48690 12936 48694 12992
rect 48694 12936 48750 12992
rect 48750 12936 48754 12992
rect 48690 12932 48754 12936
rect 48770 12992 48834 12996
rect 48770 12936 48774 12992
rect 48774 12936 48830 12992
rect 48830 12936 48834 12992
rect 48770 12932 48834 12936
rect 48850 12992 48914 12996
rect 48850 12936 48854 12992
rect 48854 12936 48910 12992
rect 48910 12936 48914 12992
rect 48850 12932 48914 12936
rect 48930 12992 48994 12996
rect 48930 12936 48934 12992
rect 48934 12936 48990 12992
rect 48990 12936 48994 12992
rect 48930 12932 48994 12936
rect 46702 12877 46766 12881
rect 46702 12821 46706 12877
rect 46706 12821 46762 12877
rect 46762 12821 46766 12877
rect 46702 12817 46766 12821
rect 46782 12877 46846 12881
rect 46782 12821 46786 12877
rect 46786 12821 46842 12877
rect 46842 12821 46846 12877
rect 46782 12817 46846 12821
rect 46862 12877 46926 12881
rect 46862 12821 46866 12877
rect 46866 12821 46922 12877
rect 46922 12821 46926 12877
rect 46862 12817 46926 12821
rect 46942 12877 47006 12881
rect 46942 12821 46946 12877
rect 46946 12821 47002 12877
rect 47002 12821 47006 12877
rect 46942 12817 47006 12821
rect 47368 12877 47432 12881
rect 47368 12821 47372 12877
rect 47372 12821 47428 12877
rect 47428 12821 47432 12877
rect 47368 12817 47432 12821
rect 47448 12877 47512 12881
rect 47448 12821 47452 12877
rect 47452 12821 47508 12877
rect 47508 12821 47512 12877
rect 47448 12817 47512 12821
rect 47528 12877 47592 12881
rect 47528 12821 47532 12877
rect 47532 12821 47588 12877
rect 47588 12821 47592 12877
rect 47528 12817 47592 12821
rect 47608 12877 47672 12881
rect 47608 12821 47612 12877
rect 47612 12821 47668 12877
rect 47668 12821 47672 12877
rect 47608 12817 47672 12821
rect 48027 12873 48091 12877
rect 48027 12817 48031 12873
rect 48031 12817 48087 12873
rect 48087 12817 48091 12873
rect 48027 12813 48091 12817
rect 48107 12873 48171 12877
rect 48107 12817 48111 12873
rect 48111 12817 48167 12873
rect 48167 12817 48171 12873
rect 48107 12813 48171 12817
rect 48187 12873 48251 12877
rect 48187 12817 48191 12873
rect 48191 12817 48247 12873
rect 48247 12817 48251 12873
rect 48187 12813 48251 12817
rect 48267 12873 48331 12877
rect 48267 12817 48271 12873
rect 48271 12817 48327 12873
rect 48327 12817 48331 12873
rect 48267 12813 48331 12817
rect 48690 12873 48754 12877
rect 48690 12817 48694 12873
rect 48694 12817 48750 12873
rect 48750 12817 48754 12873
rect 48690 12813 48754 12817
rect 48770 12873 48834 12877
rect 48770 12817 48774 12873
rect 48774 12817 48830 12873
rect 48830 12817 48834 12873
rect 48770 12813 48834 12817
rect 48850 12873 48914 12877
rect 48850 12817 48854 12873
rect 48854 12817 48910 12873
rect 48910 12817 48914 12873
rect 48850 12813 48914 12817
rect 48930 12873 48994 12877
rect 48930 12817 48934 12873
rect 48934 12817 48990 12873
rect 48990 12817 48994 12873
rect 48930 12813 48994 12817
rect 50831 13108 50895 13112
rect 50831 13052 50835 13108
rect 50835 13052 50891 13108
rect 50891 13052 50895 13108
rect 50831 13048 50895 13052
rect 50911 13108 50975 13112
rect 50911 13052 50915 13108
rect 50915 13052 50971 13108
rect 50971 13052 50975 13108
rect 50911 13048 50975 13052
rect 50991 13108 51055 13112
rect 50991 13052 50995 13108
rect 50995 13052 51051 13108
rect 51051 13052 51055 13108
rect 50991 13048 51055 13052
rect 51071 13108 51135 13112
rect 51071 13052 51075 13108
rect 51075 13052 51131 13108
rect 51131 13052 51135 13108
rect 51071 13048 51135 13052
rect 51497 13108 51561 13112
rect 51497 13052 51501 13108
rect 51501 13052 51557 13108
rect 51557 13052 51561 13108
rect 51497 13048 51561 13052
rect 51577 13108 51641 13112
rect 51577 13052 51581 13108
rect 51581 13052 51637 13108
rect 51637 13052 51641 13108
rect 51577 13048 51641 13052
rect 51657 13108 51721 13112
rect 51657 13052 51661 13108
rect 51661 13052 51717 13108
rect 51717 13052 51721 13108
rect 51657 13048 51721 13052
rect 51737 13108 51801 13112
rect 51737 13052 51741 13108
rect 51741 13052 51797 13108
rect 51797 13052 51801 13108
rect 51737 13048 51801 13052
rect 52156 13104 52220 13108
rect 52156 13048 52160 13104
rect 52160 13048 52216 13104
rect 52216 13048 52220 13104
rect 52156 13044 52220 13048
rect 52236 13104 52300 13108
rect 52236 13048 52240 13104
rect 52240 13048 52296 13104
rect 52296 13048 52300 13104
rect 52236 13044 52300 13048
rect 52316 13104 52380 13108
rect 52316 13048 52320 13104
rect 52320 13048 52376 13104
rect 52376 13048 52380 13104
rect 52316 13044 52380 13048
rect 52396 13104 52460 13108
rect 52396 13048 52400 13104
rect 52400 13048 52456 13104
rect 52456 13048 52460 13104
rect 52396 13044 52460 13048
rect 52819 13104 52883 13108
rect 52819 13048 52823 13104
rect 52823 13048 52879 13104
rect 52879 13048 52883 13104
rect 52819 13044 52883 13048
rect 52899 13104 52963 13108
rect 52899 13048 52903 13104
rect 52903 13048 52959 13104
rect 52959 13048 52963 13104
rect 52899 13044 52963 13048
rect 52979 13104 53043 13108
rect 52979 13048 52983 13104
rect 52983 13048 53039 13104
rect 53039 13048 53043 13104
rect 52979 13044 53043 13048
rect 53059 13104 53123 13108
rect 53059 13048 53063 13104
rect 53063 13048 53119 13104
rect 53119 13048 53123 13104
rect 53059 13044 53123 13048
rect 50831 12996 50895 13000
rect 50831 12940 50835 12996
rect 50835 12940 50891 12996
rect 50891 12940 50895 12996
rect 50831 12936 50895 12940
rect 50911 12996 50975 13000
rect 50911 12940 50915 12996
rect 50915 12940 50971 12996
rect 50971 12940 50975 12996
rect 50911 12936 50975 12940
rect 50991 12996 51055 13000
rect 50991 12940 50995 12996
rect 50995 12940 51051 12996
rect 51051 12940 51055 12996
rect 50991 12936 51055 12940
rect 51071 12996 51135 13000
rect 51071 12940 51075 12996
rect 51075 12940 51131 12996
rect 51131 12940 51135 12996
rect 51071 12936 51135 12940
rect 51497 12996 51561 13000
rect 51497 12940 51501 12996
rect 51501 12940 51557 12996
rect 51557 12940 51561 12996
rect 51497 12936 51561 12940
rect 51577 12996 51641 13000
rect 51577 12940 51581 12996
rect 51581 12940 51637 12996
rect 51637 12940 51641 12996
rect 51577 12936 51641 12940
rect 51657 12996 51721 13000
rect 51657 12940 51661 12996
rect 51661 12940 51717 12996
rect 51717 12940 51721 12996
rect 51657 12936 51721 12940
rect 51737 12996 51801 13000
rect 51737 12940 51741 12996
rect 51741 12940 51797 12996
rect 51797 12940 51801 12996
rect 51737 12936 51801 12940
rect 52156 12992 52220 12996
rect 52156 12936 52160 12992
rect 52160 12936 52216 12992
rect 52216 12936 52220 12992
rect 52156 12932 52220 12936
rect 52236 12992 52300 12996
rect 52236 12936 52240 12992
rect 52240 12936 52296 12992
rect 52296 12936 52300 12992
rect 52236 12932 52300 12936
rect 52316 12992 52380 12996
rect 52316 12936 52320 12992
rect 52320 12936 52376 12992
rect 52376 12936 52380 12992
rect 52316 12932 52380 12936
rect 52396 12992 52460 12996
rect 52396 12936 52400 12992
rect 52400 12936 52456 12992
rect 52456 12936 52460 12992
rect 52396 12932 52460 12936
rect 52819 12992 52883 12996
rect 52819 12936 52823 12992
rect 52823 12936 52879 12992
rect 52879 12936 52883 12992
rect 52819 12932 52883 12936
rect 52899 12992 52963 12996
rect 52899 12936 52903 12992
rect 52903 12936 52959 12992
rect 52959 12936 52963 12992
rect 52899 12932 52963 12936
rect 52979 12992 53043 12996
rect 52979 12936 52983 12992
rect 52983 12936 53039 12992
rect 53039 12936 53043 12992
rect 52979 12932 53043 12936
rect 53059 12992 53123 12996
rect 53059 12936 53063 12992
rect 53063 12936 53119 12992
rect 53119 12936 53123 12992
rect 53059 12932 53123 12936
rect 50831 12877 50895 12881
rect 50831 12821 50835 12877
rect 50835 12821 50891 12877
rect 50891 12821 50895 12877
rect 50831 12817 50895 12821
rect 50911 12877 50975 12881
rect 50911 12821 50915 12877
rect 50915 12821 50971 12877
rect 50971 12821 50975 12877
rect 50911 12817 50975 12821
rect 50991 12877 51055 12881
rect 50991 12821 50995 12877
rect 50995 12821 51051 12877
rect 51051 12821 51055 12877
rect 50991 12817 51055 12821
rect 51071 12877 51135 12881
rect 51071 12821 51075 12877
rect 51075 12821 51131 12877
rect 51131 12821 51135 12877
rect 51071 12817 51135 12821
rect 51497 12877 51561 12881
rect 51497 12821 51501 12877
rect 51501 12821 51557 12877
rect 51557 12821 51561 12877
rect 51497 12817 51561 12821
rect 51577 12877 51641 12881
rect 51577 12821 51581 12877
rect 51581 12821 51637 12877
rect 51637 12821 51641 12877
rect 51577 12817 51641 12821
rect 51657 12877 51721 12881
rect 51657 12821 51661 12877
rect 51661 12821 51717 12877
rect 51717 12821 51721 12877
rect 51657 12817 51721 12821
rect 51737 12877 51801 12881
rect 51737 12821 51741 12877
rect 51741 12821 51797 12877
rect 51797 12821 51801 12877
rect 51737 12817 51801 12821
rect 52156 12873 52220 12877
rect 52156 12817 52160 12873
rect 52160 12817 52216 12873
rect 52216 12817 52220 12873
rect 52156 12813 52220 12817
rect 52236 12873 52300 12877
rect 52236 12817 52240 12873
rect 52240 12817 52296 12873
rect 52296 12817 52300 12873
rect 52236 12813 52300 12817
rect 52316 12873 52380 12877
rect 52316 12817 52320 12873
rect 52320 12817 52376 12873
rect 52376 12817 52380 12873
rect 52316 12813 52380 12817
rect 52396 12873 52460 12877
rect 52396 12817 52400 12873
rect 52400 12817 52456 12873
rect 52456 12817 52460 12873
rect 52396 12813 52460 12817
rect 52819 12873 52883 12877
rect 52819 12817 52823 12873
rect 52823 12817 52879 12873
rect 52879 12817 52883 12873
rect 52819 12813 52883 12817
rect 52899 12873 52963 12877
rect 52899 12817 52903 12873
rect 52903 12817 52959 12873
rect 52959 12817 52963 12873
rect 52899 12813 52963 12817
rect 52979 12873 53043 12877
rect 52979 12817 52983 12873
rect 52983 12817 53039 12873
rect 53039 12817 53043 12873
rect 52979 12813 53043 12817
rect 53059 12873 53123 12877
rect 53059 12817 53063 12873
rect 53063 12817 53119 12873
rect 53119 12817 53123 12873
rect 53059 12813 53123 12817
<< metal4 >>
rect 31263 26804 31583 42360
rect 31263 26740 31265 26804
rect 31329 26740 31345 26804
rect 31409 26740 31425 26804
rect 31489 26740 31505 26804
rect 31569 26740 31583 26804
rect 31263 26692 31583 26740
rect 31263 26628 31265 26692
rect 31329 26628 31345 26692
rect 31409 26628 31425 26692
rect 31489 26628 31505 26692
rect 31569 26628 31583 26692
rect 31263 26573 31583 26628
rect 31263 26509 31265 26573
rect 31329 26509 31345 26573
rect 31409 26509 31425 26573
rect 31489 26509 31505 26573
rect 31569 26509 31583 26573
rect 31263 13112 31583 26509
rect 31263 13048 31265 13112
rect 31329 13048 31345 13112
rect 31409 13048 31425 13112
rect 31489 13048 31505 13112
rect 31569 13048 31583 13112
rect 31263 13000 31583 13048
rect 31263 12936 31265 13000
rect 31329 12936 31345 13000
rect 31409 12936 31425 13000
rect 31489 12936 31505 13000
rect 31569 12936 31583 13000
rect 31263 12881 31583 12936
rect 31263 12817 31265 12881
rect 31329 12817 31345 12881
rect 31409 12817 31425 12881
rect 31489 12817 31505 12881
rect 31569 12817 31583 12881
rect 31263 660 31583 12817
rect 31923 26804 32243 42360
rect 31923 26740 31931 26804
rect 31995 26740 32011 26804
rect 32075 26740 32091 26804
rect 32155 26740 32171 26804
rect 32235 26740 32243 26804
rect 31923 26692 32243 26740
rect 31923 26628 31931 26692
rect 31995 26628 32011 26692
rect 32075 26628 32091 26692
rect 32155 26628 32171 26692
rect 32235 26628 32243 26692
rect 31923 26573 32243 26628
rect 31923 26509 31931 26573
rect 31995 26509 32011 26573
rect 32075 26509 32091 26573
rect 32155 26509 32171 26573
rect 32235 26509 32243 26573
rect 31923 13112 32243 26509
rect 31923 13048 31931 13112
rect 31995 13048 32011 13112
rect 32075 13048 32091 13112
rect 32155 13048 32171 13112
rect 32235 13048 32243 13112
rect 31923 13000 32243 13048
rect 31923 12936 31931 13000
rect 31995 12936 32011 13000
rect 32075 12936 32091 13000
rect 32155 12936 32171 13000
rect 32235 12936 32243 13000
rect 31923 12881 32243 12936
rect 31923 12817 31931 12881
rect 31995 12817 32011 12881
rect 32075 12817 32091 12881
rect 32155 12817 32171 12881
rect 32235 12817 32243 12881
rect 31923 660 32243 12817
rect 32583 26800 32903 42360
rect 32583 26736 32590 26800
rect 32654 26736 32670 26800
rect 32734 26736 32750 26800
rect 32814 26736 32830 26800
rect 32894 26736 32903 26800
rect 32583 26688 32903 26736
rect 32583 26624 32590 26688
rect 32654 26624 32670 26688
rect 32734 26624 32750 26688
rect 32814 26624 32830 26688
rect 32894 26624 32903 26688
rect 32583 26569 32903 26624
rect 32583 26505 32590 26569
rect 32654 26505 32670 26569
rect 32734 26505 32750 26569
rect 32814 26505 32830 26569
rect 32894 26505 32903 26569
rect 32583 13108 32903 26505
rect 32583 13044 32590 13108
rect 32654 13044 32670 13108
rect 32734 13044 32750 13108
rect 32814 13044 32830 13108
rect 32894 13044 32903 13108
rect 32583 12996 32903 13044
rect 32583 12932 32590 12996
rect 32654 12932 32670 12996
rect 32734 12932 32750 12996
rect 32814 12932 32830 12996
rect 32894 12932 32903 12996
rect 32583 12877 32903 12932
rect 32583 12813 32590 12877
rect 32654 12813 32670 12877
rect 32734 12813 32750 12877
rect 32814 12813 32830 12877
rect 32894 12813 32903 12877
rect 32583 660 32903 12813
rect 33243 26800 33563 42360
rect 33243 26736 33253 26800
rect 33317 26736 33333 26800
rect 33397 26736 33413 26800
rect 33477 26736 33493 26800
rect 33557 26736 33563 26800
rect 33243 26688 33563 26736
rect 33243 26624 33253 26688
rect 33317 26624 33333 26688
rect 33397 26624 33413 26688
rect 33477 26624 33493 26688
rect 33557 26624 33563 26688
rect 33243 26569 33563 26624
rect 33243 26505 33253 26569
rect 33317 26505 33333 26569
rect 33397 26505 33413 26569
rect 33477 26505 33493 26569
rect 33557 26505 33563 26569
rect 33243 13108 33563 26505
rect 33243 13044 33253 13108
rect 33317 13044 33333 13108
rect 33397 13044 33413 13108
rect 33477 13044 33493 13108
rect 33557 13044 33563 13108
rect 33243 12996 33563 13044
rect 33243 12932 33253 12996
rect 33317 12932 33333 12996
rect 33397 12932 33413 12996
rect 33477 12932 33493 12996
rect 33557 12932 33563 12996
rect 33243 12877 33563 12932
rect 33243 12813 33253 12877
rect 33317 12813 33333 12877
rect 33397 12813 33413 12877
rect 33477 12813 33493 12877
rect 33557 12813 33563 12877
rect 33243 660 33563 12813
rect 35387 26804 35707 42360
rect 35387 26740 35394 26804
rect 35458 26740 35474 26804
rect 35538 26740 35554 26804
rect 35618 26740 35634 26804
rect 35698 26740 35707 26804
rect 35387 26692 35707 26740
rect 35387 26628 35394 26692
rect 35458 26628 35474 26692
rect 35538 26628 35554 26692
rect 35618 26628 35634 26692
rect 35698 26628 35707 26692
rect 35387 26573 35707 26628
rect 35387 26509 35394 26573
rect 35458 26509 35474 26573
rect 35538 26509 35554 26573
rect 35618 26509 35634 26573
rect 35698 26509 35707 26573
rect 35387 13112 35707 26509
rect 35387 13048 35394 13112
rect 35458 13048 35474 13112
rect 35538 13048 35554 13112
rect 35618 13048 35634 13112
rect 35698 13048 35707 13112
rect 35387 13000 35707 13048
rect 35387 12936 35394 13000
rect 35458 12936 35474 13000
rect 35538 12936 35554 13000
rect 35618 12936 35634 13000
rect 35698 12936 35707 13000
rect 35387 12881 35707 12936
rect 35387 12817 35394 12881
rect 35458 12817 35474 12881
rect 35538 12817 35554 12881
rect 35618 12817 35634 12881
rect 35698 12817 35707 12881
rect 35387 660 35707 12817
rect 36047 26804 36367 42360
rect 36047 26740 36060 26804
rect 36124 26740 36140 26804
rect 36204 26740 36220 26804
rect 36284 26740 36300 26804
rect 36364 26740 36367 26804
rect 36047 26692 36367 26740
rect 36047 26628 36060 26692
rect 36124 26628 36140 26692
rect 36204 26628 36220 26692
rect 36284 26628 36300 26692
rect 36364 26628 36367 26692
rect 36047 26573 36367 26628
rect 36047 26509 36060 26573
rect 36124 26509 36140 26573
rect 36204 26509 36220 26573
rect 36284 26509 36300 26573
rect 36364 26509 36367 26573
rect 36047 13112 36367 26509
rect 36047 13048 36060 13112
rect 36124 13048 36140 13112
rect 36204 13048 36220 13112
rect 36284 13048 36300 13112
rect 36364 13048 36367 13112
rect 36047 13000 36367 13048
rect 36047 12936 36060 13000
rect 36124 12936 36140 13000
rect 36204 12936 36220 13000
rect 36284 12936 36300 13000
rect 36364 12936 36367 13000
rect 36047 12881 36367 12936
rect 36047 12817 36060 12881
rect 36124 12817 36140 12881
rect 36204 12817 36220 12881
rect 36284 12817 36300 12881
rect 36364 12817 36367 12881
rect 36047 660 36367 12817
rect 36707 26800 37027 42360
rect 36707 26736 36719 26800
rect 36783 26736 36799 26800
rect 36863 26736 36879 26800
rect 36943 26736 36959 26800
rect 37023 26736 37027 26800
rect 36707 26688 37027 26736
rect 36707 26624 36719 26688
rect 36783 26624 36799 26688
rect 36863 26624 36879 26688
rect 36943 26624 36959 26688
rect 37023 26624 37027 26688
rect 36707 26569 37027 26624
rect 36707 26505 36719 26569
rect 36783 26505 36799 26569
rect 36863 26505 36879 26569
rect 36943 26505 36959 26569
rect 37023 26505 37027 26569
rect 36707 13108 37027 26505
rect 36707 13044 36719 13108
rect 36783 13044 36799 13108
rect 36863 13044 36879 13108
rect 36943 13044 36959 13108
rect 37023 13044 37027 13108
rect 36707 12996 37027 13044
rect 36707 12932 36719 12996
rect 36783 12932 36799 12996
rect 36863 12932 36879 12996
rect 36943 12932 36959 12996
rect 37023 12932 37027 12996
rect 36707 12877 37027 12932
rect 36707 12813 36719 12877
rect 36783 12813 36799 12877
rect 36863 12813 36879 12877
rect 36943 12813 36959 12877
rect 37023 12813 37027 12877
rect 36707 660 37027 12813
rect 37367 26800 37687 42360
rect 37367 26736 37382 26800
rect 37446 26736 37462 26800
rect 37526 26736 37542 26800
rect 37606 26736 37622 26800
rect 37686 26736 37687 26800
rect 37367 26688 37687 26736
rect 37367 26624 37382 26688
rect 37446 26624 37462 26688
rect 37526 26624 37542 26688
rect 37606 26624 37622 26688
rect 37686 26624 37687 26688
rect 37367 26569 37687 26624
rect 37367 26505 37382 26569
rect 37446 26505 37462 26569
rect 37526 26505 37542 26569
rect 37606 26505 37622 26569
rect 37686 26505 37687 26569
rect 37367 13108 37687 26505
rect 37367 13044 37382 13108
rect 37446 13044 37462 13108
rect 37526 13044 37542 13108
rect 37606 13044 37622 13108
rect 37686 13044 37687 13108
rect 37367 12996 37687 13044
rect 37367 12932 37382 12996
rect 37446 12932 37462 12996
rect 37526 12932 37542 12996
rect 37606 12932 37622 12996
rect 37686 12932 37687 12996
rect 37367 12877 37687 12932
rect 37367 12813 37382 12877
rect 37446 12813 37462 12877
rect 37526 12813 37542 12877
rect 37606 12813 37622 12877
rect 37686 12813 37687 12877
rect 37367 660 37687 12813
rect 40221 13624 40541 42360
rect 40221 13560 40315 13624
rect 40379 13560 40395 13624
rect 40459 13560 40541 13624
rect 40221 13505 40541 13560
rect 40221 13441 40315 13505
rect 40379 13441 40395 13505
rect 40459 13441 40541 13505
rect 40221 13384 40541 13441
rect 40221 13320 40315 13384
rect 40379 13320 40395 13384
rect 40459 13320 40541 13384
rect 40221 13277 40541 13320
rect 40221 13213 40315 13277
rect 40379 13213 40395 13277
rect 40459 13213 40541 13277
rect 40221 13151 40541 13213
rect 40221 13087 40315 13151
rect 40379 13087 40395 13151
rect 40459 13087 40541 13151
rect 40221 13039 40541 13087
rect 40221 12975 40315 13039
rect 40379 12975 40395 13039
rect 40459 12975 40541 13039
rect 40221 12920 40541 12975
rect 40221 12856 40315 12920
rect 40379 12856 40395 12920
rect 40459 12856 40541 12920
rect 40221 660 40541 12856
rect 42688 13568 43008 42360
rect 42688 13504 42790 13568
rect 42854 13504 42870 13568
rect 42934 13504 43008 13568
rect 42688 13445 43008 13504
rect 42688 13381 42790 13445
rect 42854 13381 42870 13445
rect 42934 13381 43008 13445
rect 42688 13333 43008 13381
rect 42688 13269 42790 13333
rect 42854 13269 42870 13333
rect 42934 13269 43008 13333
rect 42688 13214 43008 13269
rect 42688 13150 42790 13214
rect 42854 13150 42870 13214
rect 42934 13150 43008 13214
rect 42688 13090 43008 13150
rect 42688 13026 42790 13090
rect 42854 13026 42870 13090
rect 42934 13026 43008 13090
rect 42688 12983 43008 13026
rect 42688 12919 42790 12983
rect 42854 12919 42870 12983
rect 42934 12919 43008 12983
rect 42688 660 43008 12919
rect 46700 26804 47020 42360
rect 46700 26740 46702 26804
rect 46766 26740 46782 26804
rect 46846 26740 46862 26804
rect 46926 26740 46942 26804
rect 47006 26740 47020 26804
rect 46700 26692 47020 26740
rect 46700 26628 46702 26692
rect 46766 26628 46782 26692
rect 46846 26628 46862 26692
rect 46926 26628 46942 26692
rect 47006 26628 47020 26692
rect 46700 26573 47020 26628
rect 46700 26509 46702 26573
rect 46766 26509 46782 26573
rect 46846 26509 46862 26573
rect 46926 26509 46942 26573
rect 47006 26509 47020 26573
rect 46700 13112 47020 26509
rect 46700 13048 46702 13112
rect 46766 13048 46782 13112
rect 46846 13048 46862 13112
rect 46926 13048 46942 13112
rect 47006 13048 47020 13112
rect 46700 13000 47020 13048
rect 46700 12936 46702 13000
rect 46766 12936 46782 13000
rect 46846 12936 46862 13000
rect 46926 12936 46942 13000
rect 47006 12936 47020 13000
rect 46700 12881 47020 12936
rect 46700 12817 46702 12881
rect 46766 12817 46782 12881
rect 46846 12817 46862 12881
rect 46926 12817 46942 12881
rect 47006 12817 47020 12881
rect 46700 660 47020 12817
rect 47360 26804 47680 42360
rect 47360 26740 47368 26804
rect 47432 26740 47448 26804
rect 47512 26740 47528 26804
rect 47592 26740 47608 26804
rect 47672 26740 47680 26804
rect 47360 26692 47680 26740
rect 47360 26628 47368 26692
rect 47432 26628 47448 26692
rect 47512 26628 47528 26692
rect 47592 26628 47608 26692
rect 47672 26628 47680 26692
rect 47360 26573 47680 26628
rect 47360 26509 47368 26573
rect 47432 26509 47448 26573
rect 47512 26509 47528 26573
rect 47592 26509 47608 26573
rect 47672 26509 47680 26573
rect 47360 13112 47680 26509
rect 47360 13048 47368 13112
rect 47432 13048 47448 13112
rect 47512 13048 47528 13112
rect 47592 13048 47608 13112
rect 47672 13048 47680 13112
rect 47360 13000 47680 13048
rect 47360 12936 47368 13000
rect 47432 12936 47448 13000
rect 47512 12936 47528 13000
rect 47592 12936 47608 13000
rect 47672 12936 47680 13000
rect 47360 12881 47680 12936
rect 47360 12817 47368 12881
rect 47432 12817 47448 12881
rect 47512 12817 47528 12881
rect 47592 12817 47608 12881
rect 47672 12817 47680 12881
rect 47360 660 47680 12817
rect 48020 26800 48340 42360
rect 48020 26736 48027 26800
rect 48091 26736 48107 26800
rect 48171 26736 48187 26800
rect 48251 26736 48267 26800
rect 48331 26736 48340 26800
rect 48020 26688 48340 26736
rect 48020 26624 48027 26688
rect 48091 26624 48107 26688
rect 48171 26624 48187 26688
rect 48251 26624 48267 26688
rect 48331 26624 48340 26688
rect 48020 26569 48340 26624
rect 48020 26505 48027 26569
rect 48091 26505 48107 26569
rect 48171 26505 48187 26569
rect 48251 26505 48267 26569
rect 48331 26505 48340 26569
rect 48020 13108 48340 26505
rect 48020 13044 48027 13108
rect 48091 13044 48107 13108
rect 48171 13044 48187 13108
rect 48251 13044 48267 13108
rect 48331 13044 48340 13108
rect 48020 12996 48340 13044
rect 48020 12932 48027 12996
rect 48091 12932 48107 12996
rect 48171 12932 48187 12996
rect 48251 12932 48267 12996
rect 48331 12932 48340 12996
rect 48020 12877 48340 12932
rect 48020 12813 48027 12877
rect 48091 12813 48107 12877
rect 48171 12813 48187 12877
rect 48251 12813 48267 12877
rect 48331 12813 48340 12877
rect 48020 660 48340 12813
rect 48680 26800 49000 42360
rect 48680 26736 48690 26800
rect 48754 26736 48770 26800
rect 48834 26736 48850 26800
rect 48914 26736 48930 26800
rect 48994 26736 49000 26800
rect 48680 26688 49000 26736
rect 48680 26624 48690 26688
rect 48754 26624 48770 26688
rect 48834 26624 48850 26688
rect 48914 26624 48930 26688
rect 48994 26624 49000 26688
rect 48680 26569 49000 26624
rect 48680 26505 48690 26569
rect 48754 26505 48770 26569
rect 48834 26505 48850 26569
rect 48914 26505 48930 26569
rect 48994 26505 49000 26569
rect 48680 13108 49000 26505
rect 48680 13044 48690 13108
rect 48754 13044 48770 13108
rect 48834 13044 48850 13108
rect 48914 13044 48930 13108
rect 48994 13044 49000 13108
rect 48680 12996 49000 13044
rect 48680 12932 48690 12996
rect 48754 12932 48770 12996
rect 48834 12932 48850 12996
rect 48914 12932 48930 12996
rect 48994 12932 49000 12996
rect 48680 12877 49000 12932
rect 48680 12813 48690 12877
rect 48754 12813 48770 12877
rect 48834 12813 48850 12877
rect 48914 12813 48930 12877
rect 48994 12813 49000 12877
rect 48680 660 49000 12813
rect 50824 26804 51144 42360
rect 50824 26740 50831 26804
rect 50895 26740 50911 26804
rect 50975 26740 50991 26804
rect 51055 26740 51071 26804
rect 51135 26740 51144 26804
rect 50824 26692 51144 26740
rect 50824 26628 50831 26692
rect 50895 26628 50911 26692
rect 50975 26628 50991 26692
rect 51055 26628 51071 26692
rect 51135 26628 51144 26692
rect 50824 26573 51144 26628
rect 50824 26509 50831 26573
rect 50895 26509 50911 26573
rect 50975 26509 50991 26573
rect 51055 26509 51071 26573
rect 51135 26509 51144 26573
rect 50824 13112 51144 26509
rect 50824 13048 50831 13112
rect 50895 13048 50911 13112
rect 50975 13048 50991 13112
rect 51055 13048 51071 13112
rect 51135 13048 51144 13112
rect 50824 13000 51144 13048
rect 50824 12936 50831 13000
rect 50895 12936 50911 13000
rect 50975 12936 50991 13000
rect 51055 12936 51071 13000
rect 51135 12936 51144 13000
rect 50824 12881 51144 12936
rect 50824 12817 50831 12881
rect 50895 12817 50911 12881
rect 50975 12817 50991 12881
rect 51055 12817 51071 12881
rect 51135 12817 51144 12881
rect 50824 660 51144 12817
rect 51484 26804 51804 42360
rect 51484 26740 51497 26804
rect 51561 26740 51577 26804
rect 51641 26740 51657 26804
rect 51721 26740 51737 26804
rect 51801 26740 51804 26804
rect 51484 26692 51804 26740
rect 51484 26628 51497 26692
rect 51561 26628 51577 26692
rect 51641 26628 51657 26692
rect 51721 26628 51737 26692
rect 51801 26628 51804 26692
rect 51484 26573 51804 26628
rect 51484 26509 51497 26573
rect 51561 26509 51577 26573
rect 51641 26509 51657 26573
rect 51721 26509 51737 26573
rect 51801 26509 51804 26573
rect 51484 13112 51804 26509
rect 51484 13048 51497 13112
rect 51561 13048 51577 13112
rect 51641 13048 51657 13112
rect 51721 13048 51737 13112
rect 51801 13048 51804 13112
rect 51484 13000 51804 13048
rect 51484 12936 51497 13000
rect 51561 12936 51577 13000
rect 51641 12936 51657 13000
rect 51721 12936 51737 13000
rect 51801 12936 51804 13000
rect 51484 12881 51804 12936
rect 51484 12817 51497 12881
rect 51561 12817 51577 12881
rect 51641 12817 51657 12881
rect 51721 12817 51737 12881
rect 51801 12817 51804 12881
rect 51484 660 51804 12817
rect 52144 26800 52464 42360
rect 52144 26736 52156 26800
rect 52220 26736 52236 26800
rect 52300 26736 52316 26800
rect 52380 26736 52396 26800
rect 52460 26736 52464 26800
rect 52144 26688 52464 26736
rect 52144 26624 52156 26688
rect 52220 26624 52236 26688
rect 52300 26624 52316 26688
rect 52380 26624 52396 26688
rect 52460 26624 52464 26688
rect 52144 26569 52464 26624
rect 52144 26505 52156 26569
rect 52220 26505 52236 26569
rect 52300 26505 52316 26569
rect 52380 26505 52396 26569
rect 52460 26505 52464 26569
rect 52144 13108 52464 26505
rect 52144 13044 52156 13108
rect 52220 13044 52236 13108
rect 52300 13044 52316 13108
rect 52380 13044 52396 13108
rect 52460 13044 52464 13108
rect 52144 12996 52464 13044
rect 52144 12932 52156 12996
rect 52220 12932 52236 12996
rect 52300 12932 52316 12996
rect 52380 12932 52396 12996
rect 52460 12932 52464 12996
rect 52144 12877 52464 12932
rect 52144 12813 52156 12877
rect 52220 12813 52236 12877
rect 52300 12813 52316 12877
rect 52380 12813 52396 12877
rect 52460 12813 52464 12877
rect 52144 660 52464 12813
rect 52804 26800 53124 42360
rect 52804 26736 52819 26800
rect 52883 26736 52899 26800
rect 52963 26736 52979 26800
rect 53043 26736 53059 26800
rect 53123 26736 53124 26800
rect 52804 26688 53124 26736
rect 52804 26624 52819 26688
rect 52883 26624 52899 26688
rect 52963 26624 52979 26688
rect 53043 26624 53059 26688
rect 53123 26624 53124 26688
rect 52804 26569 53124 26624
rect 52804 26505 52819 26569
rect 52883 26505 52899 26569
rect 52963 26505 52979 26569
rect 53043 26505 53059 26569
rect 53123 26505 53124 26569
rect 52804 13108 53124 26505
rect 52804 13044 52819 13108
rect 52883 13044 52899 13108
rect 52963 13044 52979 13108
rect 53043 13044 53059 13108
rect 53123 13044 53124 13108
rect 52804 12996 53124 13044
rect 52804 12932 52819 12996
rect 52883 12932 52899 12996
rect 52963 12932 52979 12996
rect 53043 12932 53059 12996
rect 53123 12932 53124 12996
rect 52804 12877 53124 12932
rect 52804 12813 52819 12877
rect 52883 12813 52899 12877
rect 52963 12813 52979 12877
rect 53043 12813 53059 12877
rect 53123 12813 53124 12877
rect 52804 660 53124 12813
use sky130_ef_ip__xtal_osc_32k  mprj
timestamp 1527873355
transform 0 -1 67059 -1 0 26820
box 0 11646 14034 38204
<< labels >>
flabel metal2 s 1365 42249 1493 43705 0 FreeSans 280 90 0 0 in
port 4 nsew
flabel metal2 s 103165 42249 103293 43705 0 FreeSans 280 90 0 0 out
port 3 nsew
flabel metal2 s 43239 -656 43295 144 0 FreeSans 280 90 0 0 boost
port 1 nsew
flabel metal2 s 40756 -656 40812 144 0 FreeSans 280 90 0 0 ena
port 2 nsew
flabel metal2 s 39916 -656 39972 144 0 FreeSans 280 90 0 0 dout
port 5 nsew
flabel metal4 s 33243 660 33563 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 31923 660 32243 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 31263 660 31583 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 32583 660 32903 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 37367 660 37687 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 36047 660 36367 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 35387 660 35707 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 36707 660 37027 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 48680 660 49000 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 47360 660 47680 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 48020 660 48340 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
flabel metal4 s 51484 660 51804 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 50824 660 51144 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 52144 660 52464 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 40221 660 40541 42360 0 FreeSans 2400 90 0 0 vssd1
port 8 nsew
flabel metal4 s 42688 660 43008 42360 0 FreeSans 2400 90 0 0 vccd1
port 9 nsew
flabel metal4 s 52804 660 53124 42360 0 FreeSans 2400 90 0 0 vdda1
port 6 nsew
flabel metal4 s 46700 660 47020 42360 0 FreeSans 2400 90 0 0 vssa1
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 105060 42360
<< end >>
