VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_32k_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_32k_DI ;
  ORIGIN -58.230 0.000 ;
  SIZE 525.300 BY 211.800 ;
  PIN boost
    ANTENNAGATEAREA 0.510000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 277.560 75.500 277.730 76.000 ;
        RECT 278.530 75.500 278.700 76.000 ;
        RECT 278.585 71.080 278.915 71.570 ;
        RECT 274.055 67.310 274.225 67.640 ;
        RECT 275.650 67.310 275.820 67.640 ;
      LAYER mcon ;
        RECT 277.560 75.665 277.730 75.835 ;
        RECT 278.530 75.665 278.700 75.835 ;
        RECT 278.665 71.240 278.835 71.410 ;
        RECT 274.055 67.390 274.225 67.560 ;
        RECT 275.650 67.390 275.820 67.560 ;
      LAYER met1 ;
        RECT 275.620 75.820 275.950 75.870 ;
        RECT 277.530 75.820 277.760 75.980 ;
        RECT 278.500 75.820 278.730 75.980 ;
        RECT 275.620 75.620 278.730 75.820 ;
        RECT 275.620 75.280 275.950 75.620 ;
        RECT 277.520 75.520 277.760 75.620 ;
        RECT 278.500 75.520 278.730 75.620 ;
        RECT 275.705 71.480 275.975 71.845 ;
        RECT 278.555 71.480 278.945 71.550 ;
        RECT 275.705 71.220 278.945 71.480 ;
        RECT 275.705 71.170 275.975 71.220 ;
        RECT 278.555 71.100 278.945 71.220 ;
        RECT 274.025 67.550 274.255 67.620 ;
        RECT 274.670 67.550 275.040 67.600 ;
        RECT 275.620 67.550 275.850 67.620 ;
        RECT 274.010 67.310 275.870 67.550 ;
        RECT 274.670 67.130 275.040 67.310 ;
        RECT 274.360 66.130 275.360 67.130 ;
      LAYER via ;
        RECT 275.655 75.445 275.915 75.705 ;
        RECT 275.710 71.380 275.970 71.640 ;
        RECT 274.725 67.220 274.985 67.480 ;
      LAYER met2 ;
        RECT 275.570 75.330 276.000 75.820 ;
        RECT 275.660 71.795 275.930 75.330 ;
        RECT 275.655 71.220 276.025 71.795 ;
        RECT 275.660 68.490 275.930 71.220 ;
        RECT 274.725 68.220 275.930 68.490 ;
        RECT 274.725 67.865 274.995 68.220 ;
        RECT 274.725 67.550 275.040 67.865 ;
        RECT 274.620 67.150 275.090 67.550 ;
        RECT 274.770 64.930 275.040 67.150 ;
        RECT 274.425 0.000 275.425 64.930 ;
        RECT 274.425 -3.280 274.705 0.000 ;
    END
  END boost
  PIN ena
    ANTENNAGATEAREA 0.585000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 259.340 75.500 259.510 76.000 ;
        RECT 260.310 75.500 260.480 76.000 ;
        RECT 262.220 67.310 262.390 67.640 ;
        RECT 263.815 67.310 263.985 67.640 ;
        RECT 261.210 64.930 261.540 65.420 ;
        RECT 267.885 64.820 268.055 65.150 ;
      LAYER mcon ;
        RECT 259.340 75.665 259.510 75.835 ;
        RECT 260.310 75.665 260.480 75.835 ;
        RECT 262.220 67.390 262.390 67.560 ;
        RECT 263.815 67.390 263.985 67.560 ;
        RECT 261.290 65.090 261.460 65.260 ;
        RECT 267.885 64.900 268.055 65.070 ;
      LAYER met1 ;
        RECT 259.310 75.820 259.540 75.980 ;
        RECT 260.280 75.820 260.510 75.980 ;
        RECT 262.090 75.820 262.420 75.870 ;
        RECT 259.310 75.620 262.420 75.820 ;
        RECT 259.310 75.520 259.540 75.620 ;
        RECT 260.280 75.520 260.520 75.620 ;
        RECT 262.090 75.280 262.420 75.620 ;
        RECT 262.190 67.550 262.420 67.620 ;
        RECT 263.000 67.550 263.370 67.600 ;
        RECT 263.785 67.550 264.015 67.620 ;
        RECT 262.170 67.310 264.030 67.550 ;
        RECT 263.000 67.130 263.370 67.310 ;
        RECT 262.680 66.130 263.680 67.130 ;
        RECT 262.680 66.120 262.965 66.130 ;
        RECT 261.290 65.875 262.965 66.120 ;
        RECT 261.290 65.400 261.535 65.875 ;
        RECT 262.680 65.800 262.965 65.875 ;
        RECT 267.800 65.790 268.060 66.150 ;
        RECT 261.180 64.950 261.570 65.400 ;
        RECT 267.860 65.130 268.060 65.790 ;
        RECT 267.855 64.840 268.085 65.130 ;
      LAYER via ;
        RECT 262.125 75.445 262.385 75.705 ;
        RECT 263.055 67.220 263.315 67.480 ;
        RECT 262.695 65.875 262.955 66.135 ;
        RECT 267.800 65.840 268.060 66.100 ;
      LAYER met2 ;
        RECT 262.040 75.330 262.470 75.820 ;
        RECT 262.110 68.490 262.380 75.330 ;
        RECT 262.110 68.220 263.315 68.490 ;
        RECT 263.045 67.550 263.315 68.220 ;
        RECT 262.950 67.150 263.420 67.550 ;
        RECT 262.630 66.100 263.015 66.150 ;
        RECT 262.630 65.905 268.150 66.100 ;
        RECT 262.630 65.855 263.015 65.905 ;
        RECT 262.680 64.930 262.965 65.855 ;
        RECT 267.750 65.840 268.110 65.905 ;
        RECT 262.010 0.000 263.010 64.930 ;
        RECT 262.010 -3.280 262.290 0.000 ;
    END
  END ena
  PIN out
    PORT
      LAYER met2 ;
        RECT 574.055 166.965 574.695 218.525 ;
        RECT 279.250 165.865 574.695 166.965 ;
        RECT 279.250 133.100 280.250 165.865 ;
    END
  END out
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER li1 ;
        RECT 270.115 90.280 270.285 90.780 ;
        RECT 276.775 90.040 277.235 90.210 ;
        RECT 266.840 88.900 267.010 89.400 ;
        RECT 257.780 88.055 258.110 88.545 ;
        RECT 205.335 84.500 207.495 84.850 ;
        RECT 257.765 84.785 258.095 85.275 ;
      LAYER mcon ;
        RECT 270.115 90.445 270.285 90.615 ;
        RECT 276.920 90.040 277.090 90.210 ;
        RECT 266.840 89.065 267.010 89.235 ;
        RECT 257.860 88.215 258.030 88.385 ;
        RECT 257.845 84.945 258.015 85.115 ;
        RECT 205.435 84.590 205.605 84.760 ;
        RECT 205.795 84.590 205.965 84.760 ;
        RECT 206.155 84.590 206.325 84.760 ;
        RECT 206.515 84.590 206.685 84.760 ;
        RECT 206.875 84.590 207.045 84.760 ;
        RECT 207.235 84.590 207.405 84.760 ;
      LAYER met1 ;
        RECT 203.400 133.100 204.400 134.100 ;
        RECT 203.655 83.415 204.090 133.100 ;
        RECT 270.085 90.590 270.315 90.760 ;
        RECT 268.390 90.385 270.315 90.590 ;
        RECT 266.810 89.250 267.040 89.380 ;
        RECT 268.390 89.250 268.595 90.385 ;
        RECT 270.085 90.300 270.315 90.385 ;
        RECT 276.795 90.010 277.215 90.240 ;
        RECT 266.810 89.235 268.595 89.250 ;
        RECT 272.620 89.235 273.505 89.340 ;
        RECT 266.810 89.045 273.505 89.235 ;
        RECT 266.810 88.920 267.040 89.045 ;
        RECT 268.335 89.030 273.505 89.045 ;
        RECT 257.765 88.525 258.110 88.565 ;
        RECT 257.750 88.075 258.140 88.525 ;
        RECT 257.765 85.255 258.110 88.075 ;
        RECT 268.335 87.700 268.650 89.030 ;
        RECT 272.620 88.885 273.505 89.030 ;
        RECT 274.875 89.280 275.760 89.335 ;
        RECT 276.855 89.280 277.095 90.010 ;
        RECT 274.875 89.040 277.095 89.280 ;
        RECT 274.875 88.880 275.760 89.040 ;
        RECT 268.345 85.360 268.660 86.575 ;
        RECT 205.335 83.415 207.495 84.850 ;
        RECT 257.735 84.805 258.125 85.255 ;
        RECT 257.765 83.415 258.110 84.805 ;
        RECT 268.370 84.345 268.640 85.360 ;
        RECT 203.655 83.385 258.110 83.415 ;
        RECT 263.440 84.075 268.640 84.345 ;
        RECT 263.440 83.385 263.710 84.075 ;
        RECT 203.655 83.115 263.710 83.385 ;
        RECT 203.655 83.030 258.110 83.115 ;
        RECT 203.655 82.980 258.105 83.030 ;
      LAYER via ;
        RECT 203.615 133.325 204.195 133.905 ;
        RECT 272.775 88.985 273.035 89.245 ;
        RECT 273.095 88.985 273.355 89.245 ;
        RECT 275.030 88.980 275.290 89.240 ;
        RECT 275.350 88.980 275.610 89.240 ;
        RECT 268.365 88.500 268.625 88.760 ;
        RECT 268.365 88.180 268.625 88.440 ;
        RECT 268.365 87.860 268.625 88.120 ;
        RECT 268.375 86.160 268.635 86.420 ;
        RECT 268.375 85.840 268.635 86.100 ;
        RECT 268.375 85.520 268.635 85.780 ;
      LAYER met2 ;
        RECT 65.055 142.320 65.695 218.525 ;
        RECT 65.055 141.080 204.400 142.320 ;
        RECT 203.400 133.100 204.400 141.080 ;
        POLYGON 204.400 142.320 204.405 142.320 204.400 133.905 ;
        RECT 272.570 89.245 273.555 89.290 ;
        RECT 274.825 89.245 275.810 89.285 ;
        RECT 272.570 89.005 275.810 89.245 ;
        RECT 272.570 88.935 273.555 89.005 ;
        RECT 274.825 88.930 275.810 89.005 ;
        RECT 268.285 87.750 268.700 88.865 ;
        RECT 268.305 86.525 268.680 87.750 ;
        RECT 268.295 85.410 268.710 86.525 ;
    END
  END in
  PIN dout
    PORT
      LAYER li1 ;
        RECT 262.025 70.320 264.185 71.010 ;
      LAYER mcon ;
        RECT 262.120 70.400 264.090 70.930 ;
      LAYER met1 ;
        RECT 262.055 70.865 264.160 70.960 ;
        RECT 258.085 70.480 264.160 70.865 ;
        RECT 258.085 64.930 258.470 70.480 ;
        RECT 262.055 70.370 264.160 70.480 ;
        RECT 257.810 63.930 258.810 64.930 ;
      LAYER via ;
        RECT 258.005 64.155 258.585 64.735 ;
      LAYER met2 ;
        RECT 257.810 0.000 258.810 64.930 ;
        RECT 257.810 -3.280 258.090 0.000 ;
    END
  END dout
  PIN vdda1
    ANTENNADIFFAREA 200.228592 ;
    PORT
      LAYER nwell ;
        RECT 202.505 132.520 335.295 134.100 ;
        RECT 202.505 65.510 204.085 132.520 ;
        RECT 257.015 84.115 258.845 85.945 ;
        RECT 261.665 84.070 268.095 99.930 ;
        RECT 261.720 77.250 276.320 80.330 ;
        RECT 261.730 74.060 276.310 77.250 ;
        RECT 255.535 72.480 282.295 74.060 ;
        RECT 255.535 65.510 257.115 72.480 ;
        RECT 202.505 63.930 257.115 65.510 ;
        RECT 280.715 65.510 282.295 72.480 ;
        RECT 333.565 65.510 335.295 132.520 ;
        RECT 280.715 63.930 335.295 65.510 ;
      LAYER li1 ;
        RECT 209.405 133.665 229.825 133.815 ;
        RECT 230.855 133.665 250.675 133.770 ;
        RECT 251.410 133.665 278.040 133.815 ;
        RECT 308.095 133.665 328.000 133.765 ;
        RECT 330.225 133.665 332.375 133.770 ;
        RECT 202.940 133.495 334.860 133.665 ;
        RECT 202.940 130.945 203.110 133.495 ;
        RECT 209.405 133.395 229.825 133.495 ;
        RECT 230.855 133.395 250.675 133.495 ;
        RECT 251.410 133.380 278.040 133.495 ;
        RECT 308.095 133.390 328.000 133.495 ;
        RECT 330.225 133.395 332.375 133.495 ;
        RECT 334.690 133.225 334.860 133.495 ;
        RECT 330.225 131.200 332.385 131.550 ;
        RECT 202.835 65.265 203.165 130.945 ;
        RECT 267.595 99.540 268.200 99.560 ;
        RECT 265.445 99.505 268.200 99.540 ;
        RECT 261.250 99.370 268.200 99.505 ;
        RECT 261.250 97.410 265.615 99.370 ;
        RECT 267.535 97.410 268.200 99.370 ;
        RECT 261.250 96.290 268.200 97.410 ;
        RECT 261.250 94.330 262.225 96.290 ;
        RECT 263.135 95.620 263.595 95.790 ;
        RECT 264.145 94.330 265.615 96.290 ;
        RECT 267.535 94.330 268.200 96.290 ;
        RECT 261.250 93.210 268.200 94.330 ;
        RECT 261.250 91.250 262.225 93.210 ;
        RECT 263.135 92.540 263.595 92.710 ;
        RECT 264.145 91.250 265.615 93.210 ;
        RECT 267.535 91.250 268.200 93.210 ;
        RECT 261.250 90.130 268.200 91.250 ;
        RECT 261.250 88.170 262.225 90.130 ;
        RECT 263.135 89.460 263.595 89.630 ;
        RECT 264.145 88.170 265.615 90.130 ;
        RECT 267.535 88.170 268.200 90.130 ;
        RECT 261.250 87.050 268.200 88.170 ;
        RECT 257.195 85.760 258.665 85.765 ;
        RECT 257.195 85.595 258.905 85.760 ;
        RECT 257.195 84.465 257.365 85.595 ;
        RECT 258.495 84.465 258.905 85.595 ;
        RECT 257.195 84.295 258.905 84.465 ;
        RECT 261.250 85.090 262.225 87.050 ;
        RECT 263.135 85.590 263.595 85.760 ;
        RECT 264.145 85.090 265.615 87.050 ;
        RECT 266.165 85.590 266.625 85.760 ;
        RECT 267.535 85.090 268.200 87.050 ;
        RECT 261.250 84.420 268.200 85.090 ;
        RECT 258.495 84.290 258.905 84.295 ;
        RECT 261.760 79.730 268.510 80.360 ;
        RECT 261.760 77.810 262.300 79.730 ;
        RECT 264.550 77.810 265.630 79.730 ;
        RECT 266.535 78.310 266.995 78.480 ;
        RECT 267.890 77.810 268.510 79.730 ;
        RECT 261.760 76.720 268.510 77.810 ;
        RECT 261.760 74.760 262.300 76.720 ;
        RECT 264.560 76.690 268.510 76.720 ;
        RECT 264.560 74.760 265.630 76.690 ;
        RECT 266.535 76.020 266.995 76.190 ;
        RECT 261.760 74.750 265.630 74.760 ;
        RECT 267.890 74.750 268.510 76.690 ;
        RECT 261.760 74.120 268.510 74.750 ;
        RECT 269.530 79.730 276.280 80.360 ;
        RECT 269.530 77.810 270.150 79.730 ;
        RECT 271.045 78.310 271.505 78.480 ;
        RECT 272.410 77.810 273.490 79.730 ;
        RECT 275.740 77.810 276.280 79.730 ;
        RECT 269.530 76.720 276.280 77.810 ;
        RECT 269.530 76.690 273.480 76.720 ;
        RECT 269.530 74.750 270.150 76.690 ;
        RECT 271.045 76.020 271.505 76.190 ;
        RECT 272.410 74.760 273.480 76.690 ;
        RECT 275.740 74.760 276.280 76.720 ;
        RECT 272.410 74.750 276.280 74.760 ;
        RECT 269.530 74.120 276.280 74.750 ;
        RECT 256.940 73.135 280.975 73.200 ;
        RECT 256.500 72.965 281.380 73.135 ;
        RECT 256.500 72.235 256.670 72.965 ;
        RECT 256.940 72.900 280.975 72.965 ;
        RECT 281.210 72.395 281.380 72.965 ;
        RECT 205.385 66.560 207.545 66.910 ;
        RECT 202.940 64.535 203.110 65.265 ;
        RECT 256.415 64.905 256.735 72.235 ;
        RECT 281.115 65.210 281.405 72.395 ;
        RECT 205.385 64.535 207.540 64.640 ;
        RECT 209.365 64.535 229.275 64.625 ;
        RECT 230.875 64.535 250.705 64.635 ;
        RECT 251.455 64.535 256.110 64.645 ;
        RECT 256.500 64.535 256.670 64.905 ;
        RECT 202.940 64.365 256.670 64.535 ;
        RECT 281.210 64.535 281.380 65.210 ;
        RECT 334.575 64.835 334.955 133.225 ;
        RECT 282.080 64.535 306.415 64.665 ;
        RECT 308.155 64.535 327.985 64.630 ;
        RECT 334.690 64.535 334.860 64.835 ;
        RECT 281.210 64.365 334.860 64.535 ;
        RECT 205.385 64.265 207.540 64.365 ;
        RECT 209.365 64.255 229.275 64.365 ;
        RECT 230.875 64.265 250.705 64.365 ;
        RECT 251.455 64.270 256.110 64.365 ;
        RECT 282.080 64.350 306.415 64.365 ;
        RECT 308.155 64.265 327.985 64.365 ;
      LAYER mcon ;
        RECT 209.450 133.520 209.620 133.690 ;
        RECT 209.810 133.520 209.980 133.690 ;
        RECT 210.170 133.520 210.340 133.690 ;
        RECT 210.530 133.520 210.700 133.690 ;
        RECT 210.890 133.520 211.060 133.690 ;
        RECT 211.250 133.520 211.420 133.690 ;
        RECT 211.610 133.520 211.780 133.690 ;
        RECT 211.970 133.520 212.140 133.690 ;
        RECT 212.330 133.520 212.500 133.690 ;
        RECT 212.690 133.520 212.860 133.690 ;
        RECT 213.050 133.520 213.220 133.690 ;
        RECT 213.410 133.520 213.580 133.690 ;
        RECT 213.770 133.520 213.940 133.690 ;
        RECT 214.130 133.520 214.300 133.690 ;
        RECT 214.490 133.520 214.660 133.690 ;
        RECT 214.850 133.520 215.020 133.690 ;
        RECT 215.210 133.520 215.380 133.690 ;
        RECT 215.570 133.520 215.740 133.690 ;
        RECT 215.930 133.520 216.100 133.690 ;
        RECT 216.290 133.520 216.460 133.690 ;
        RECT 216.650 133.520 216.820 133.690 ;
        RECT 217.010 133.520 217.180 133.690 ;
        RECT 217.370 133.520 217.540 133.690 ;
        RECT 217.730 133.520 217.900 133.690 ;
        RECT 218.090 133.520 218.260 133.690 ;
        RECT 218.450 133.520 218.620 133.690 ;
        RECT 218.810 133.520 218.980 133.690 ;
        RECT 219.170 133.520 219.340 133.690 ;
        RECT 219.530 133.520 219.700 133.690 ;
        RECT 219.890 133.520 220.060 133.690 ;
        RECT 220.250 133.520 220.420 133.690 ;
        RECT 220.610 133.520 220.780 133.690 ;
        RECT 220.970 133.520 221.140 133.690 ;
        RECT 221.330 133.520 221.500 133.690 ;
        RECT 221.690 133.520 221.860 133.690 ;
        RECT 222.050 133.520 222.220 133.690 ;
        RECT 222.410 133.520 222.580 133.690 ;
        RECT 222.770 133.520 222.940 133.690 ;
        RECT 223.130 133.520 223.300 133.690 ;
        RECT 223.490 133.520 223.660 133.690 ;
        RECT 223.850 133.520 224.020 133.690 ;
        RECT 224.210 133.520 224.380 133.690 ;
        RECT 224.570 133.520 224.740 133.690 ;
        RECT 224.930 133.520 225.100 133.690 ;
        RECT 225.290 133.520 225.460 133.690 ;
        RECT 225.650 133.520 225.820 133.690 ;
        RECT 226.010 133.520 226.180 133.690 ;
        RECT 226.370 133.520 226.540 133.690 ;
        RECT 226.730 133.520 226.900 133.690 ;
        RECT 227.090 133.520 227.260 133.690 ;
        RECT 227.450 133.520 227.620 133.690 ;
        RECT 227.810 133.520 227.980 133.690 ;
        RECT 228.170 133.520 228.340 133.690 ;
        RECT 228.530 133.520 228.700 133.690 ;
        RECT 228.890 133.520 229.060 133.690 ;
        RECT 229.250 133.520 229.420 133.690 ;
        RECT 229.610 133.520 229.780 133.690 ;
        RECT 230.960 133.500 231.130 133.670 ;
        RECT 231.320 133.500 231.490 133.670 ;
        RECT 231.680 133.500 231.850 133.670 ;
        RECT 232.040 133.500 232.210 133.670 ;
        RECT 232.400 133.500 232.570 133.670 ;
        RECT 232.760 133.500 232.930 133.670 ;
        RECT 233.120 133.500 233.290 133.670 ;
        RECT 233.480 133.500 233.650 133.670 ;
        RECT 233.840 133.500 234.010 133.670 ;
        RECT 234.200 133.500 234.370 133.670 ;
        RECT 234.560 133.500 234.730 133.670 ;
        RECT 234.920 133.500 235.090 133.670 ;
        RECT 235.280 133.500 235.450 133.670 ;
        RECT 235.640 133.500 235.810 133.670 ;
        RECT 236.000 133.500 236.170 133.670 ;
        RECT 236.360 133.500 236.530 133.670 ;
        RECT 236.720 133.500 236.890 133.670 ;
        RECT 237.080 133.500 237.250 133.670 ;
        RECT 237.440 133.500 237.610 133.670 ;
        RECT 237.800 133.500 237.970 133.670 ;
        RECT 238.160 133.500 238.330 133.670 ;
        RECT 238.520 133.500 238.690 133.670 ;
        RECT 238.880 133.500 239.050 133.670 ;
        RECT 239.240 133.500 239.410 133.670 ;
        RECT 239.600 133.500 239.770 133.670 ;
        RECT 239.960 133.500 240.130 133.670 ;
        RECT 240.320 133.500 240.490 133.670 ;
        RECT 240.680 133.500 240.850 133.670 ;
        RECT 241.040 133.500 241.210 133.670 ;
        RECT 241.400 133.500 241.570 133.670 ;
        RECT 241.760 133.500 241.930 133.670 ;
        RECT 242.120 133.500 242.290 133.670 ;
        RECT 242.480 133.500 242.650 133.670 ;
        RECT 242.840 133.500 243.010 133.670 ;
        RECT 243.200 133.500 243.370 133.670 ;
        RECT 243.560 133.500 243.730 133.670 ;
        RECT 243.920 133.500 244.090 133.670 ;
        RECT 244.280 133.500 244.450 133.670 ;
        RECT 244.640 133.500 244.810 133.670 ;
        RECT 245.000 133.500 245.170 133.670 ;
        RECT 245.360 133.500 245.530 133.670 ;
        RECT 245.720 133.500 245.890 133.670 ;
        RECT 246.080 133.500 246.250 133.670 ;
        RECT 246.440 133.500 246.610 133.670 ;
        RECT 246.800 133.500 246.970 133.670 ;
        RECT 247.160 133.500 247.330 133.670 ;
        RECT 247.520 133.500 247.690 133.670 ;
        RECT 247.880 133.500 248.050 133.670 ;
        RECT 248.240 133.500 248.410 133.670 ;
        RECT 248.600 133.500 248.770 133.670 ;
        RECT 248.960 133.500 249.130 133.670 ;
        RECT 249.320 133.500 249.490 133.670 ;
        RECT 249.680 133.500 249.850 133.670 ;
        RECT 250.040 133.500 250.210 133.670 ;
        RECT 250.400 133.500 250.570 133.670 ;
        RECT 251.500 133.515 251.670 133.685 ;
        RECT 251.860 133.515 252.030 133.685 ;
        RECT 252.220 133.515 252.390 133.685 ;
        RECT 252.580 133.515 252.750 133.685 ;
        RECT 252.940 133.515 253.110 133.685 ;
        RECT 253.300 133.515 253.470 133.685 ;
        RECT 253.660 133.515 253.830 133.685 ;
        RECT 254.020 133.515 254.190 133.685 ;
        RECT 254.380 133.515 254.550 133.685 ;
        RECT 254.740 133.515 254.910 133.685 ;
        RECT 255.100 133.515 255.270 133.685 ;
        RECT 255.460 133.515 255.630 133.685 ;
        RECT 255.820 133.515 255.990 133.685 ;
        RECT 256.180 133.515 256.350 133.685 ;
        RECT 256.540 133.515 256.710 133.685 ;
        RECT 256.900 133.515 257.070 133.685 ;
        RECT 257.260 133.515 257.430 133.685 ;
        RECT 257.620 133.515 257.790 133.685 ;
        RECT 257.980 133.515 258.150 133.685 ;
        RECT 258.340 133.515 258.510 133.685 ;
        RECT 258.700 133.515 258.870 133.685 ;
        RECT 259.060 133.515 259.230 133.685 ;
        RECT 259.420 133.515 259.590 133.685 ;
        RECT 259.780 133.515 259.950 133.685 ;
        RECT 260.140 133.515 260.310 133.685 ;
        RECT 260.500 133.515 260.670 133.685 ;
        RECT 260.860 133.515 261.030 133.685 ;
        RECT 261.220 133.515 261.390 133.685 ;
        RECT 261.580 133.515 261.750 133.685 ;
        RECT 261.940 133.515 262.110 133.685 ;
        RECT 262.300 133.515 262.470 133.685 ;
        RECT 262.660 133.515 262.830 133.685 ;
        RECT 263.020 133.515 263.190 133.685 ;
        RECT 263.380 133.515 263.550 133.685 ;
        RECT 263.740 133.515 263.910 133.685 ;
        RECT 264.100 133.515 264.270 133.685 ;
        RECT 264.460 133.515 264.630 133.685 ;
        RECT 264.820 133.515 264.990 133.685 ;
        RECT 265.180 133.515 265.350 133.685 ;
        RECT 265.540 133.515 265.710 133.685 ;
        RECT 265.900 133.515 266.070 133.685 ;
        RECT 266.260 133.515 266.430 133.685 ;
        RECT 266.620 133.515 266.790 133.685 ;
        RECT 266.980 133.515 267.150 133.685 ;
        RECT 267.340 133.515 267.510 133.685 ;
        RECT 267.700 133.515 267.870 133.685 ;
        RECT 268.060 133.515 268.230 133.685 ;
        RECT 268.420 133.515 268.590 133.685 ;
        RECT 268.780 133.515 268.950 133.685 ;
        RECT 269.140 133.515 269.310 133.685 ;
        RECT 269.500 133.515 269.670 133.685 ;
        RECT 269.860 133.515 270.030 133.685 ;
        RECT 270.220 133.515 270.390 133.685 ;
        RECT 270.580 133.515 270.750 133.685 ;
        RECT 270.940 133.515 271.110 133.685 ;
        RECT 271.300 133.515 271.470 133.685 ;
        RECT 271.660 133.515 271.830 133.685 ;
        RECT 272.020 133.515 272.190 133.685 ;
        RECT 272.380 133.515 272.550 133.685 ;
        RECT 272.740 133.515 272.910 133.685 ;
        RECT 273.100 133.515 273.270 133.685 ;
        RECT 273.460 133.515 273.630 133.685 ;
        RECT 273.820 133.515 273.990 133.685 ;
        RECT 274.180 133.515 274.350 133.685 ;
        RECT 274.540 133.515 274.710 133.685 ;
        RECT 274.900 133.515 275.070 133.685 ;
        RECT 275.260 133.515 275.430 133.685 ;
        RECT 275.620 133.515 275.790 133.685 ;
        RECT 275.980 133.515 276.150 133.685 ;
        RECT 276.340 133.515 276.510 133.685 ;
        RECT 276.700 133.515 276.870 133.685 ;
        RECT 277.060 133.515 277.230 133.685 ;
        RECT 277.420 133.515 277.590 133.685 ;
        RECT 277.780 133.515 277.950 133.685 ;
        RECT 308.245 133.495 308.415 133.665 ;
        RECT 308.605 133.495 308.775 133.665 ;
        RECT 308.965 133.495 309.135 133.665 ;
        RECT 309.325 133.495 309.495 133.665 ;
        RECT 309.685 133.495 309.855 133.665 ;
        RECT 310.045 133.495 310.215 133.665 ;
        RECT 310.405 133.495 310.575 133.665 ;
        RECT 310.765 133.495 310.935 133.665 ;
        RECT 311.125 133.495 311.295 133.665 ;
        RECT 311.485 133.495 311.655 133.665 ;
        RECT 311.845 133.495 312.015 133.665 ;
        RECT 312.205 133.495 312.375 133.665 ;
        RECT 312.565 133.495 312.735 133.665 ;
        RECT 312.925 133.495 313.095 133.665 ;
        RECT 313.285 133.495 313.455 133.665 ;
        RECT 313.645 133.495 313.815 133.665 ;
        RECT 314.005 133.495 314.175 133.665 ;
        RECT 314.365 133.495 314.535 133.665 ;
        RECT 314.725 133.495 314.895 133.665 ;
        RECT 315.085 133.495 315.255 133.665 ;
        RECT 315.445 133.495 315.615 133.665 ;
        RECT 315.805 133.495 315.975 133.665 ;
        RECT 316.165 133.495 316.335 133.665 ;
        RECT 316.525 133.495 316.695 133.665 ;
        RECT 316.885 133.495 317.055 133.665 ;
        RECT 317.245 133.495 317.415 133.665 ;
        RECT 317.605 133.495 317.775 133.665 ;
        RECT 317.965 133.495 318.135 133.665 ;
        RECT 318.325 133.495 318.495 133.665 ;
        RECT 318.685 133.495 318.855 133.665 ;
        RECT 319.045 133.495 319.215 133.665 ;
        RECT 319.405 133.495 319.575 133.665 ;
        RECT 319.765 133.495 319.935 133.665 ;
        RECT 320.125 133.495 320.295 133.665 ;
        RECT 320.485 133.495 320.655 133.665 ;
        RECT 320.845 133.495 321.015 133.665 ;
        RECT 321.205 133.495 321.375 133.665 ;
        RECT 321.565 133.495 321.735 133.665 ;
        RECT 321.925 133.495 322.095 133.665 ;
        RECT 322.285 133.495 322.455 133.665 ;
        RECT 322.645 133.495 322.815 133.665 ;
        RECT 323.005 133.495 323.175 133.665 ;
        RECT 323.365 133.495 323.535 133.665 ;
        RECT 323.725 133.495 323.895 133.665 ;
        RECT 324.085 133.495 324.255 133.665 ;
        RECT 324.445 133.495 324.615 133.665 ;
        RECT 324.805 133.495 324.975 133.665 ;
        RECT 325.165 133.495 325.335 133.665 ;
        RECT 325.525 133.495 325.695 133.665 ;
        RECT 325.885 133.495 326.055 133.665 ;
        RECT 326.245 133.495 326.415 133.665 ;
        RECT 326.605 133.495 326.775 133.665 ;
        RECT 326.965 133.495 327.135 133.665 ;
        RECT 327.325 133.495 327.495 133.665 ;
        RECT 327.685 133.495 327.855 133.665 ;
        RECT 330.315 133.500 330.485 133.670 ;
        RECT 330.675 133.500 330.845 133.670 ;
        RECT 331.035 133.500 331.205 133.670 ;
        RECT 331.395 133.500 331.565 133.670 ;
        RECT 331.755 133.500 331.925 133.670 ;
        RECT 332.115 133.500 332.285 133.670 ;
        RECT 334.680 132.965 334.850 133.135 ;
        RECT 334.680 132.605 334.850 132.775 ;
        RECT 334.680 132.245 334.850 132.415 ;
        RECT 334.680 131.885 334.850 132.055 ;
        RECT 330.320 131.290 330.490 131.460 ;
        RECT 330.680 131.290 330.850 131.460 ;
        RECT 331.040 131.290 331.210 131.460 ;
        RECT 331.400 131.290 331.570 131.460 ;
        RECT 331.760 131.290 331.930 131.460 ;
        RECT 332.120 131.290 332.290 131.460 ;
        RECT 334.680 131.525 334.850 131.695 ;
        RECT 334.680 131.165 334.850 131.335 ;
        RECT 202.915 130.600 203.085 130.770 ;
        RECT 202.915 130.240 203.085 130.410 ;
        RECT 202.915 129.880 203.085 130.050 ;
        RECT 202.915 129.520 203.085 129.690 ;
        RECT 202.915 129.160 203.085 129.330 ;
        RECT 202.915 128.800 203.085 128.970 ;
        RECT 202.915 128.440 203.085 128.610 ;
        RECT 202.915 128.080 203.085 128.250 ;
        RECT 202.915 127.720 203.085 127.890 ;
        RECT 202.915 127.360 203.085 127.530 ;
        RECT 202.915 127.000 203.085 127.170 ;
        RECT 202.915 126.640 203.085 126.810 ;
        RECT 202.915 126.280 203.085 126.450 ;
        RECT 202.915 125.920 203.085 126.090 ;
        RECT 202.915 125.560 203.085 125.730 ;
        RECT 202.915 125.200 203.085 125.370 ;
        RECT 202.915 124.840 203.085 125.010 ;
        RECT 202.915 124.480 203.085 124.650 ;
        RECT 202.915 124.120 203.085 124.290 ;
        RECT 202.915 123.760 203.085 123.930 ;
        RECT 202.915 123.400 203.085 123.570 ;
        RECT 202.915 123.040 203.085 123.210 ;
        RECT 202.915 122.680 203.085 122.850 ;
        RECT 202.915 122.320 203.085 122.490 ;
        RECT 202.915 121.960 203.085 122.130 ;
        RECT 202.915 121.600 203.085 121.770 ;
        RECT 202.915 121.240 203.085 121.410 ;
        RECT 202.915 120.880 203.085 121.050 ;
        RECT 202.915 120.520 203.085 120.690 ;
        RECT 202.915 120.160 203.085 120.330 ;
        RECT 202.915 119.800 203.085 119.970 ;
        RECT 202.915 119.440 203.085 119.610 ;
        RECT 202.915 119.080 203.085 119.250 ;
        RECT 202.915 118.720 203.085 118.890 ;
        RECT 202.915 118.360 203.085 118.530 ;
        RECT 202.915 118.000 203.085 118.170 ;
        RECT 202.915 117.640 203.085 117.810 ;
        RECT 202.915 117.280 203.085 117.450 ;
        RECT 202.915 116.920 203.085 117.090 ;
        RECT 202.915 116.560 203.085 116.730 ;
        RECT 202.915 116.200 203.085 116.370 ;
        RECT 202.915 115.840 203.085 116.010 ;
        RECT 202.915 115.480 203.085 115.650 ;
        RECT 202.915 115.120 203.085 115.290 ;
        RECT 202.915 114.760 203.085 114.930 ;
        RECT 202.915 114.400 203.085 114.570 ;
        RECT 202.915 114.040 203.085 114.210 ;
        RECT 202.915 113.680 203.085 113.850 ;
        RECT 202.915 113.320 203.085 113.490 ;
        RECT 202.915 112.960 203.085 113.130 ;
        RECT 202.915 112.600 203.085 112.770 ;
        RECT 202.915 112.240 203.085 112.410 ;
        RECT 202.915 111.880 203.085 112.050 ;
        RECT 202.915 111.520 203.085 111.690 ;
        RECT 202.915 111.160 203.085 111.330 ;
        RECT 202.915 110.800 203.085 110.970 ;
        RECT 202.915 110.440 203.085 110.610 ;
        RECT 202.915 110.080 203.085 110.250 ;
        RECT 202.915 109.720 203.085 109.890 ;
        RECT 202.915 109.360 203.085 109.530 ;
        RECT 202.915 109.000 203.085 109.170 ;
        RECT 202.915 108.640 203.085 108.810 ;
        RECT 202.915 108.280 203.085 108.450 ;
        RECT 202.915 107.920 203.085 108.090 ;
        RECT 202.915 107.560 203.085 107.730 ;
        RECT 202.915 107.200 203.085 107.370 ;
        RECT 202.915 106.840 203.085 107.010 ;
        RECT 202.915 106.480 203.085 106.650 ;
        RECT 202.915 106.120 203.085 106.290 ;
        RECT 202.915 105.760 203.085 105.930 ;
        RECT 202.915 105.400 203.085 105.570 ;
        RECT 202.915 105.040 203.085 105.210 ;
        RECT 202.915 104.680 203.085 104.850 ;
        RECT 202.915 104.320 203.085 104.490 ;
        RECT 202.915 103.960 203.085 104.130 ;
        RECT 202.915 103.600 203.085 103.770 ;
        RECT 202.915 103.240 203.085 103.410 ;
        RECT 202.915 102.880 203.085 103.050 ;
        RECT 202.915 102.520 203.085 102.690 ;
        RECT 202.915 102.160 203.085 102.330 ;
        RECT 202.915 101.800 203.085 101.970 ;
        RECT 202.915 101.440 203.085 101.610 ;
        RECT 202.915 101.080 203.085 101.250 ;
        RECT 202.915 100.720 203.085 100.890 ;
        RECT 202.915 100.360 203.085 100.530 ;
        RECT 202.915 100.000 203.085 100.170 ;
        RECT 202.915 99.640 203.085 99.810 ;
        RECT 334.680 130.805 334.850 130.975 ;
        RECT 334.680 130.445 334.850 130.615 ;
        RECT 334.680 130.085 334.850 130.255 ;
        RECT 334.680 129.725 334.850 129.895 ;
        RECT 334.680 129.365 334.850 129.535 ;
        RECT 334.680 129.005 334.850 129.175 ;
        RECT 334.680 128.645 334.850 128.815 ;
        RECT 334.680 128.285 334.850 128.455 ;
        RECT 334.680 127.925 334.850 128.095 ;
        RECT 334.680 127.565 334.850 127.735 ;
        RECT 334.680 127.205 334.850 127.375 ;
        RECT 334.680 126.845 334.850 127.015 ;
        RECT 334.680 126.485 334.850 126.655 ;
        RECT 334.680 126.125 334.850 126.295 ;
        RECT 334.680 125.765 334.850 125.935 ;
        RECT 334.680 125.405 334.850 125.575 ;
        RECT 334.680 125.045 334.850 125.215 ;
        RECT 334.680 124.685 334.850 124.855 ;
        RECT 334.680 124.325 334.850 124.495 ;
        RECT 334.680 123.965 334.850 124.135 ;
        RECT 334.680 123.605 334.850 123.775 ;
        RECT 334.680 123.245 334.850 123.415 ;
        RECT 334.680 122.885 334.850 123.055 ;
        RECT 334.680 122.525 334.850 122.695 ;
        RECT 334.680 122.165 334.850 122.335 ;
        RECT 334.680 121.805 334.850 121.975 ;
        RECT 334.680 121.445 334.850 121.615 ;
        RECT 334.680 121.085 334.850 121.255 ;
        RECT 334.680 120.725 334.850 120.895 ;
        RECT 334.680 120.365 334.850 120.535 ;
        RECT 334.680 120.005 334.850 120.175 ;
        RECT 334.680 119.645 334.850 119.815 ;
        RECT 334.680 119.285 334.850 119.455 ;
        RECT 334.680 118.925 334.850 119.095 ;
        RECT 334.680 118.565 334.850 118.735 ;
        RECT 334.680 118.205 334.850 118.375 ;
        RECT 334.680 117.845 334.850 118.015 ;
        RECT 334.680 117.485 334.850 117.655 ;
        RECT 334.680 117.125 334.850 117.295 ;
        RECT 334.680 116.765 334.850 116.935 ;
        RECT 334.680 116.405 334.850 116.575 ;
        RECT 334.680 116.045 334.850 116.215 ;
        RECT 334.680 115.685 334.850 115.855 ;
        RECT 334.680 115.325 334.850 115.495 ;
        RECT 334.680 114.965 334.850 115.135 ;
        RECT 334.680 114.605 334.850 114.775 ;
        RECT 334.680 114.245 334.850 114.415 ;
        RECT 334.680 113.885 334.850 114.055 ;
        RECT 334.680 113.525 334.850 113.695 ;
        RECT 334.680 113.165 334.850 113.335 ;
        RECT 334.680 112.805 334.850 112.975 ;
        RECT 334.680 112.445 334.850 112.615 ;
        RECT 334.680 112.085 334.850 112.255 ;
        RECT 334.680 111.725 334.850 111.895 ;
        RECT 334.680 111.365 334.850 111.535 ;
        RECT 334.680 111.005 334.850 111.175 ;
        RECT 334.680 110.645 334.850 110.815 ;
        RECT 334.680 110.285 334.850 110.455 ;
        RECT 334.680 109.925 334.850 110.095 ;
        RECT 334.680 109.565 334.850 109.735 ;
        RECT 334.680 109.205 334.850 109.375 ;
        RECT 334.680 108.845 334.850 109.015 ;
        RECT 334.680 108.485 334.850 108.655 ;
        RECT 334.680 108.125 334.850 108.295 ;
        RECT 334.680 107.765 334.850 107.935 ;
        RECT 334.680 107.405 334.850 107.575 ;
        RECT 334.680 107.045 334.850 107.215 ;
        RECT 334.680 106.685 334.850 106.855 ;
        RECT 334.680 106.325 334.850 106.495 ;
        RECT 334.680 105.965 334.850 106.135 ;
        RECT 334.680 105.605 334.850 105.775 ;
        RECT 334.680 105.245 334.850 105.415 ;
        RECT 334.680 104.885 334.850 105.055 ;
        RECT 334.680 104.525 334.850 104.695 ;
        RECT 334.680 104.165 334.850 104.335 ;
        RECT 334.680 103.805 334.850 103.975 ;
        RECT 334.680 103.445 334.850 103.615 ;
        RECT 334.680 103.085 334.850 103.255 ;
        RECT 334.680 102.725 334.850 102.895 ;
        RECT 334.680 102.365 334.850 102.535 ;
        RECT 334.680 102.005 334.850 102.175 ;
        RECT 334.680 101.645 334.850 101.815 ;
        RECT 334.680 101.285 334.850 101.455 ;
        RECT 334.680 100.925 334.850 101.095 ;
        RECT 334.680 100.565 334.850 100.735 ;
        RECT 334.680 100.205 334.850 100.375 ;
        RECT 334.680 99.845 334.850 100.015 ;
        RECT 202.915 99.280 203.085 99.450 ;
        RECT 202.915 98.920 203.085 99.090 ;
        RECT 202.915 98.560 203.085 98.730 ;
        RECT 202.915 98.200 203.085 98.370 ;
        RECT 202.915 97.840 203.085 98.010 ;
        RECT 202.915 97.480 203.085 97.650 ;
        RECT 202.915 97.120 203.085 97.290 ;
        RECT 202.915 96.760 203.085 96.930 ;
        RECT 202.915 96.400 203.085 96.570 ;
        RECT 202.915 96.040 203.085 96.210 ;
        RECT 202.915 95.680 203.085 95.850 ;
        RECT 202.915 95.320 203.085 95.490 ;
        RECT 202.915 94.960 203.085 95.130 ;
        RECT 202.915 94.600 203.085 94.770 ;
        RECT 202.915 94.240 203.085 94.410 ;
        RECT 202.915 93.880 203.085 94.050 ;
        RECT 202.915 93.520 203.085 93.690 ;
        RECT 202.915 93.160 203.085 93.330 ;
        RECT 202.915 92.800 203.085 92.970 ;
        RECT 202.915 92.440 203.085 92.610 ;
        RECT 202.915 92.080 203.085 92.250 ;
        RECT 202.915 91.720 203.085 91.890 ;
        RECT 202.915 91.360 203.085 91.530 ;
        RECT 202.915 91.000 203.085 91.170 ;
        RECT 202.915 90.640 203.085 90.810 ;
        RECT 202.915 90.280 203.085 90.450 ;
        RECT 202.915 89.920 203.085 90.090 ;
        RECT 202.915 89.560 203.085 89.730 ;
        RECT 202.915 89.200 203.085 89.370 ;
        RECT 202.915 88.840 203.085 89.010 ;
        RECT 202.915 88.480 203.085 88.650 ;
        RECT 202.915 88.120 203.085 88.290 ;
        RECT 202.915 87.760 203.085 87.930 ;
        RECT 202.915 87.400 203.085 87.570 ;
        RECT 202.915 87.040 203.085 87.210 ;
        RECT 202.915 86.680 203.085 86.850 ;
        RECT 202.915 86.320 203.085 86.490 ;
        RECT 202.915 85.960 203.085 86.130 ;
        RECT 202.915 85.600 203.085 85.770 ;
        RECT 264.425 98.955 264.595 99.125 ;
        RECT 264.425 98.595 264.595 98.765 ;
        RECT 264.425 98.235 264.595 98.405 ;
        RECT 264.425 97.875 264.595 98.045 ;
        RECT 264.425 97.515 264.595 97.685 ;
        RECT 264.425 97.155 264.595 97.325 ;
        RECT 264.425 96.795 264.595 96.965 ;
        RECT 263.280 95.620 263.450 95.790 ;
        RECT 264.425 95.765 264.595 95.935 ;
        RECT 264.785 95.765 264.955 95.935 ;
        RECT 265.145 95.765 265.315 95.935 ;
        RECT 263.280 92.540 263.450 92.710 ;
        RECT 264.420 92.560 264.590 92.730 ;
        RECT 264.780 92.560 264.950 92.730 ;
        RECT 265.140 92.560 265.310 92.730 ;
        RECT 263.280 89.460 263.450 89.630 ;
        RECT 264.425 89.555 264.595 89.725 ;
        RECT 264.785 89.555 264.955 89.725 ;
        RECT 265.145 89.555 265.315 89.725 ;
        RECT 202.915 85.240 203.085 85.410 ;
        RECT 202.915 84.880 203.085 85.050 ;
        RECT 202.915 84.520 203.085 84.690 ;
        RECT 202.915 84.160 203.085 84.330 ;
        RECT 258.615 85.480 258.785 85.650 ;
        RECT 258.615 85.120 258.785 85.290 ;
        RECT 258.615 84.760 258.785 84.930 ;
        RECT 258.615 84.400 258.785 84.570 ;
        RECT 263.280 85.590 263.450 85.760 ;
        RECT 266.310 85.590 266.480 85.760 ;
        RECT 264.435 85.415 264.605 85.585 ;
        RECT 264.795 85.415 264.965 85.585 ;
        RECT 265.155 85.415 265.325 85.585 ;
        RECT 334.680 99.485 334.850 99.655 ;
        RECT 334.680 99.125 334.850 99.295 ;
        RECT 334.680 98.765 334.850 98.935 ;
        RECT 334.680 98.405 334.850 98.575 ;
        RECT 334.680 98.045 334.850 98.215 ;
        RECT 334.680 97.685 334.850 97.855 ;
        RECT 334.680 97.325 334.850 97.495 ;
        RECT 334.680 96.965 334.850 97.135 ;
        RECT 334.680 96.605 334.850 96.775 ;
        RECT 334.680 96.245 334.850 96.415 ;
        RECT 334.680 95.885 334.850 96.055 ;
        RECT 334.680 95.525 334.850 95.695 ;
        RECT 334.680 95.165 334.850 95.335 ;
        RECT 334.680 94.805 334.850 94.975 ;
        RECT 334.680 94.445 334.850 94.615 ;
        RECT 334.680 94.085 334.850 94.255 ;
        RECT 334.680 93.725 334.850 93.895 ;
        RECT 334.680 93.365 334.850 93.535 ;
        RECT 334.680 93.005 334.850 93.175 ;
        RECT 334.680 92.645 334.850 92.815 ;
        RECT 334.680 92.285 334.850 92.455 ;
        RECT 334.680 91.925 334.850 92.095 ;
        RECT 334.680 91.565 334.850 91.735 ;
        RECT 334.680 91.205 334.850 91.375 ;
        RECT 334.680 90.845 334.850 91.015 ;
        RECT 334.680 90.485 334.850 90.655 ;
        RECT 334.680 90.125 334.850 90.295 ;
        RECT 334.680 89.765 334.850 89.935 ;
        RECT 334.680 89.405 334.850 89.575 ;
        RECT 334.680 89.045 334.850 89.215 ;
        RECT 334.680 88.685 334.850 88.855 ;
        RECT 334.680 88.325 334.850 88.495 ;
        RECT 334.680 87.965 334.850 88.135 ;
        RECT 334.680 87.605 334.850 87.775 ;
        RECT 334.680 87.245 334.850 87.415 ;
        RECT 334.680 86.885 334.850 87.055 ;
        RECT 334.680 86.525 334.850 86.695 ;
        RECT 334.680 86.165 334.850 86.335 ;
        RECT 334.680 85.805 334.850 85.975 ;
        RECT 334.680 85.445 334.850 85.615 ;
        RECT 334.680 85.085 334.850 85.255 ;
        RECT 334.680 84.725 334.850 84.895 ;
        RECT 334.680 84.365 334.850 84.535 ;
        RECT 202.915 83.800 203.085 83.970 ;
        RECT 202.915 83.440 203.085 83.610 ;
        RECT 202.915 83.080 203.085 83.250 ;
        RECT 202.915 82.720 203.085 82.890 ;
        RECT 202.915 82.360 203.085 82.530 ;
        RECT 202.915 82.000 203.085 82.170 ;
        RECT 202.915 81.640 203.085 81.810 ;
        RECT 202.915 81.280 203.085 81.450 ;
        RECT 202.915 80.920 203.085 81.090 ;
        RECT 202.915 80.560 203.085 80.730 ;
        RECT 202.915 80.200 203.085 80.370 ;
        RECT 334.680 84.005 334.850 84.175 ;
        RECT 334.680 83.645 334.850 83.815 ;
        RECT 334.680 83.285 334.850 83.455 ;
        RECT 334.680 82.925 334.850 83.095 ;
        RECT 334.680 82.565 334.850 82.735 ;
        RECT 334.680 82.205 334.850 82.375 ;
        RECT 334.680 81.845 334.850 82.015 ;
        RECT 334.680 81.485 334.850 81.655 ;
        RECT 334.680 81.125 334.850 81.295 ;
        RECT 334.680 80.765 334.850 80.935 ;
        RECT 334.680 80.405 334.850 80.575 ;
        RECT 202.915 79.840 203.085 80.010 ;
        RECT 202.915 79.480 203.085 79.650 ;
        RECT 202.915 79.120 203.085 79.290 ;
        RECT 202.915 78.760 203.085 78.930 ;
        RECT 202.915 78.400 203.085 78.570 ;
        RECT 202.915 78.040 203.085 78.210 ;
        RECT 202.915 77.680 203.085 77.850 ;
        RECT 202.915 77.320 203.085 77.490 ;
        RECT 202.915 76.960 203.085 77.130 ;
        RECT 202.915 76.600 203.085 76.770 ;
        RECT 202.915 76.240 203.085 76.410 ;
        RECT 202.915 75.880 203.085 76.050 ;
        RECT 202.915 75.520 203.085 75.690 ;
        RECT 202.915 75.160 203.085 75.330 ;
        RECT 202.915 74.800 203.085 74.970 ;
        RECT 202.915 74.440 203.085 74.610 ;
        RECT 202.915 74.080 203.085 74.250 ;
        RECT 267.400 79.970 267.570 80.140 ;
        RECT 267.760 79.970 267.930 80.140 ;
        RECT 268.120 79.970 268.290 80.140 ;
        RECT 266.680 78.310 266.850 78.480 ;
        RECT 266.730 76.975 268.340 77.505 ;
        RECT 266.680 76.020 266.850 76.190 ;
        RECT 267.455 74.340 267.625 74.510 ;
        RECT 267.815 74.340 267.985 74.510 ;
        RECT 268.175 74.340 268.345 74.510 ;
        RECT 269.750 79.970 269.920 80.140 ;
        RECT 270.110 79.970 270.280 80.140 ;
        RECT 270.470 79.970 270.640 80.140 ;
        RECT 271.190 78.310 271.360 78.480 ;
        RECT 269.700 76.975 271.310 77.505 ;
        RECT 271.190 76.020 271.360 76.190 ;
        RECT 269.695 74.340 269.865 74.510 ;
        RECT 270.055 74.340 270.225 74.510 ;
        RECT 270.415 74.340 270.585 74.510 ;
        RECT 334.680 80.045 334.850 80.215 ;
        RECT 334.680 79.685 334.850 79.855 ;
        RECT 334.680 79.325 334.850 79.495 ;
        RECT 334.680 78.965 334.850 79.135 ;
        RECT 334.680 78.605 334.850 78.775 ;
        RECT 334.680 78.245 334.850 78.415 ;
        RECT 334.680 77.885 334.850 78.055 ;
        RECT 334.680 77.525 334.850 77.695 ;
        RECT 334.680 77.165 334.850 77.335 ;
        RECT 334.680 76.805 334.850 76.975 ;
        RECT 334.680 76.445 334.850 76.615 ;
        RECT 334.680 76.085 334.850 76.255 ;
        RECT 334.680 75.725 334.850 75.895 ;
        RECT 334.680 75.365 334.850 75.535 ;
        RECT 334.680 75.005 334.850 75.175 ;
        RECT 334.680 74.645 334.850 74.815 ;
        RECT 334.680 74.285 334.850 74.455 ;
        RECT 202.915 73.720 203.085 73.890 ;
        RECT 202.915 73.360 203.085 73.530 ;
        RECT 334.680 73.925 334.850 74.095 ;
        RECT 334.680 73.565 334.850 73.735 ;
        RECT 334.680 73.205 334.850 73.375 ;
        RECT 202.915 73.000 203.085 73.170 ;
        RECT 202.915 72.640 203.085 72.810 ;
        RECT 202.915 72.280 203.085 72.450 ;
        RECT 256.995 72.965 257.165 73.135 ;
        RECT 257.355 72.965 257.525 73.135 ;
        RECT 257.715 72.965 257.885 73.135 ;
        RECT 258.075 72.965 258.245 73.135 ;
        RECT 258.435 72.965 258.605 73.135 ;
        RECT 258.795 72.965 258.965 73.135 ;
        RECT 259.155 72.965 259.325 73.135 ;
        RECT 259.515 72.965 259.685 73.135 ;
        RECT 259.875 72.965 260.045 73.135 ;
        RECT 260.235 72.965 260.405 73.135 ;
        RECT 260.595 72.965 260.765 73.135 ;
        RECT 260.955 72.965 261.125 73.135 ;
        RECT 261.315 72.965 261.485 73.135 ;
        RECT 261.675 72.965 261.845 73.135 ;
        RECT 262.035 72.965 262.205 73.135 ;
        RECT 262.395 72.965 262.565 73.135 ;
        RECT 262.755 72.965 262.925 73.135 ;
        RECT 263.115 72.965 263.285 73.135 ;
        RECT 263.475 72.965 263.645 73.135 ;
        RECT 263.835 72.965 264.005 73.135 ;
        RECT 264.195 72.965 264.365 73.135 ;
        RECT 264.555 72.965 264.725 73.135 ;
        RECT 264.915 72.965 265.085 73.135 ;
        RECT 265.275 72.965 265.445 73.135 ;
        RECT 265.635 72.965 265.805 73.135 ;
        RECT 265.995 72.965 266.165 73.135 ;
        RECT 266.355 72.965 266.525 73.135 ;
        RECT 266.715 72.965 266.885 73.135 ;
        RECT 267.075 72.965 267.245 73.135 ;
        RECT 267.435 72.965 267.605 73.135 ;
        RECT 267.795 72.965 267.965 73.135 ;
        RECT 268.155 72.965 268.325 73.135 ;
        RECT 268.515 72.965 268.685 73.135 ;
        RECT 268.875 72.965 269.045 73.135 ;
        RECT 269.235 72.965 269.405 73.135 ;
        RECT 269.595 72.965 269.765 73.135 ;
        RECT 269.955 72.965 270.125 73.135 ;
        RECT 270.315 72.965 270.485 73.135 ;
        RECT 270.675 72.965 270.845 73.135 ;
        RECT 271.035 72.965 271.205 73.135 ;
        RECT 271.395 72.965 271.565 73.135 ;
        RECT 271.755 72.965 271.925 73.135 ;
        RECT 272.115 72.965 272.285 73.135 ;
        RECT 272.475 72.965 272.645 73.135 ;
        RECT 272.835 72.965 273.005 73.135 ;
        RECT 273.195 72.965 273.365 73.135 ;
        RECT 273.555 72.965 273.725 73.135 ;
        RECT 273.915 72.965 274.085 73.135 ;
        RECT 274.275 72.965 274.445 73.135 ;
        RECT 274.635 72.965 274.805 73.135 ;
        RECT 274.995 72.965 275.165 73.135 ;
        RECT 275.355 72.965 275.525 73.135 ;
        RECT 275.715 72.965 275.885 73.135 ;
        RECT 276.075 72.965 276.245 73.135 ;
        RECT 276.435 72.965 276.605 73.135 ;
        RECT 276.795 72.965 276.965 73.135 ;
        RECT 277.155 72.965 277.325 73.135 ;
        RECT 277.515 72.965 277.685 73.135 ;
        RECT 277.875 72.965 278.045 73.135 ;
        RECT 278.235 72.965 278.405 73.135 ;
        RECT 278.595 72.965 278.765 73.135 ;
        RECT 278.955 72.965 279.125 73.135 ;
        RECT 279.315 72.965 279.485 73.135 ;
        RECT 279.675 72.965 279.845 73.135 ;
        RECT 280.035 72.965 280.205 73.135 ;
        RECT 280.395 72.965 280.565 73.135 ;
        RECT 280.755 72.965 280.925 73.135 ;
        RECT 334.680 72.845 334.850 73.015 ;
        RECT 334.680 72.485 334.850 72.655 ;
        RECT 202.915 71.920 203.085 72.090 ;
        RECT 202.915 71.560 203.085 71.730 ;
        RECT 202.915 71.200 203.085 71.370 ;
        RECT 202.915 70.840 203.085 71.010 ;
        RECT 202.915 70.480 203.085 70.650 ;
        RECT 202.915 70.120 203.085 70.290 ;
        RECT 202.915 69.760 203.085 69.930 ;
        RECT 202.915 69.400 203.085 69.570 ;
        RECT 202.915 69.040 203.085 69.210 ;
        RECT 202.915 68.680 203.085 68.850 ;
        RECT 202.915 68.320 203.085 68.490 ;
        RECT 202.915 67.960 203.085 68.130 ;
        RECT 202.915 67.600 203.085 67.770 ;
        RECT 202.915 67.240 203.085 67.410 ;
        RECT 202.915 66.880 203.085 67.050 ;
        RECT 256.490 71.905 256.660 72.075 ;
        RECT 256.490 71.545 256.660 71.715 ;
        RECT 256.490 71.185 256.660 71.355 ;
        RECT 256.490 70.825 256.660 70.995 ;
        RECT 256.490 70.465 256.660 70.635 ;
        RECT 256.490 70.105 256.660 70.275 ;
        RECT 256.490 69.745 256.660 69.915 ;
        RECT 256.490 69.385 256.660 69.555 ;
        RECT 256.490 69.025 256.660 69.195 ;
        RECT 256.490 68.665 256.660 68.835 ;
        RECT 256.490 68.305 256.660 68.475 ;
        RECT 256.490 67.945 256.660 68.115 ;
        RECT 256.490 67.585 256.660 67.755 ;
        RECT 256.490 67.225 256.660 67.395 ;
        RECT 202.915 66.520 203.085 66.690 ;
        RECT 205.485 66.650 205.655 66.820 ;
        RECT 205.845 66.650 206.015 66.820 ;
        RECT 206.205 66.650 206.375 66.820 ;
        RECT 206.565 66.650 206.735 66.820 ;
        RECT 206.925 66.650 207.095 66.820 ;
        RECT 207.285 66.650 207.455 66.820 ;
        RECT 256.490 66.865 256.660 67.035 ;
        RECT 202.915 66.160 203.085 66.330 ;
        RECT 202.915 65.800 203.085 65.970 ;
        RECT 202.915 65.440 203.085 65.610 ;
        RECT 256.490 66.505 256.660 66.675 ;
        RECT 256.490 66.145 256.660 66.315 ;
        RECT 256.490 65.785 256.660 65.955 ;
        RECT 256.490 65.425 256.660 65.595 ;
        RECT 256.490 65.065 256.660 65.235 ;
        RECT 281.175 72.140 281.345 72.310 ;
        RECT 281.175 71.780 281.345 71.950 ;
        RECT 281.175 71.420 281.345 71.590 ;
        RECT 281.175 71.060 281.345 71.230 ;
        RECT 281.175 70.700 281.345 70.870 ;
        RECT 281.175 70.340 281.345 70.510 ;
        RECT 281.175 69.980 281.345 70.150 ;
        RECT 281.175 69.620 281.345 69.790 ;
        RECT 281.175 69.260 281.345 69.430 ;
        RECT 281.175 68.900 281.345 69.070 ;
        RECT 281.175 68.540 281.345 68.710 ;
        RECT 281.175 68.180 281.345 68.350 ;
        RECT 281.175 67.820 281.345 67.990 ;
        RECT 281.175 67.460 281.345 67.630 ;
        RECT 281.175 67.100 281.345 67.270 ;
        RECT 281.175 66.740 281.345 66.910 ;
        RECT 281.175 66.380 281.345 66.550 ;
        RECT 281.175 66.020 281.345 66.190 ;
        RECT 281.175 65.660 281.345 65.830 ;
        RECT 281.175 65.300 281.345 65.470 ;
        RECT 334.680 72.125 334.850 72.295 ;
        RECT 334.680 71.765 334.850 71.935 ;
        RECT 334.680 71.405 334.850 71.575 ;
        RECT 334.680 71.045 334.850 71.215 ;
        RECT 334.680 70.685 334.850 70.855 ;
        RECT 334.680 70.325 334.850 70.495 ;
        RECT 334.680 69.965 334.850 70.135 ;
        RECT 334.680 69.605 334.850 69.775 ;
        RECT 334.680 69.245 334.850 69.415 ;
        RECT 334.680 68.885 334.850 69.055 ;
        RECT 334.680 68.525 334.850 68.695 ;
        RECT 334.680 68.165 334.850 68.335 ;
        RECT 334.680 67.805 334.850 67.975 ;
        RECT 334.680 67.445 334.850 67.615 ;
        RECT 334.680 67.085 334.850 67.255 ;
        RECT 334.680 66.725 334.850 66.895 ;
        RECT 334.680 66.365 334.850 66.535 ;
        RECT 334.680 66.005 334.850 66.175 ;
        RECT 334.680 65.645 334.850 65.815 ;
        RECT 334.680 65.285 334.850 65.455 ;
        RECT 205.480 64.370 205.650 64.540 ;
        RECT 205.840 64.370 206.010 64.540 ;
        RECT 206.200 64.370 206.370 64.540 ;
        RECT 206.560 64.370 206.730 64.540 ;
        RECT 206.920 64.370 207.090 64.540 ;
        RECT 207.280 64.370 207.450 64.540 ;
        RECT 209.515 64.355 209.685 64.525 ;
        RECT 209.875 64.355 210.045 64.525 ;
        RECT 210.235 64.355 210.405 64.525 ;
        RECT 210.595 64.355 210.765 64.525 ;
        RECT 210.955 64.355 211.125 64.525 ;
        RECT 211.315 64.355 211.485 64.525 ;
        RECT 211.675 64.355 211.845 64.525 ;
        RECT 212.035 64.355 212.205 64.525 ;
        RECT 212.395 64.355 212.565 64.525 ;
        RECT 212.755 64.355 212.925 64.525 ;
        RECT 213.115 64.355 213.285 64.525 ;
        RECT 213.475 64.355 213.645 64.525 ;
        RECT 213.835 64.355 214.005 64.525 ;
        RECT 214.195 64.355 214.365 64.525 ;
        RECT 214.555 64.355 214.725 64.525 ;
        RECT 214.915 64.355 215.085 64.525 ;
        RECT 215.275 64.355 215.445 64.525 ;
        RECT 215.635 64.355 215.805 64.525 ;
        RECT 215.995 64.355 216.165 64.525 ;
        RECT 216.355 64.355 216.525 64.525 ;
        RECT 216.715 64.355 216.885 64.525 ;
        RECT 217.075 64.355 217.245 64.525 ;
        RECT 217.435 64.355 217.605 64.525 ;
        RECT 217.795 64.355 217.965 64.525 ;
        RECT 218.155 64.355 218.325 64.525 ;
        RECT 218.515 64.355 218.685 64.525 ;
        RECT 218.875 64.355 219.045 64.525 ;
        RECT 219.235 64.355 219.405 64.525 ;
        RECT 219.595 64.355 219.765 64.525 ;
        RECT 219.955 64.355 220.125 64.525 ;
        RECT 220.315 64.355 220.485 64.525 ;
        RECT 220.675 64.355 220.845 64.525 ;
        RECT 221.035 64.355 221.205 64.525 ;
        RECT 221.395 64.355 221.565 64.525 ;
        RECT 221.755 64.355 221.925 64.525 ;
        RECT 222.115 64.355 222.285 64.525 ;
        RECT 222.475 64.355 222.645 64.525 ;
        RECT 222.835 64.355 223.005 64.525 ;
        RECT 223.195 64.355 223.365 64.525 ;
        RECT 223.555 64.355 223.725 64.525 ;
        RECT 223.915 64.355 224.085 64.525 ;
        RECT 224.275 64.355 224.445 64.525 ;
        RECT 224.635 64.355 224.805 64.525 ;
        RECT 224.995 64.355 225.165 64.525 ;
        RECT 225.355 64.355 225.525 64.525 ;
        RECT 225.715 64.355 225.885 64.525 ;
        RECT 226.075 64.355 226.245 64.525 ;
        RECT 226.435 64.355 226.605 64.525 ;
        RECT 226.795 64.355 226.965 64.525 ;
        RECT 227.155 64.355 227.325 64.525 ;
        RECT 227.515 64.355 227.685 64.525 ;
        RECT 227.875 64.355 228.045 64.525 ;
        RECT 228.235 64.355 228.405 64.525 ;
        RECT 228.595 64.355 228.765 64.525 ;
        RECT 228.955 64.355 229.125 64.525 ;
        RECT 230.985 64.365 231.155 64.535 ;
        RECT 231.345 64.365 231.515 64.535 ;
        RECT 231.705 64.365 231.875 64.535 ;
        RECT 232.065 64.365 232.235 64.535 ;
        RECT 232.425 64.365 232.595 64.535 ;
        RECT 232.785 64.365 232.955 64.535 ;
        RECT 233.145 64.365 233.315 64.535 ;
        RECT 233.505 64.365 233.675 64.535 ;
        RECT 233.865 64.365 234.035 64.535 ;
        RECT 234.225 64.365 234.395 64.535 ;
        RECT 234.585 64.365 234.755 64.535 ;
        RECT 234.945 64.365 235.115 64.535 ;
        RECT 235.305 64.365 235.475 64.535 ;
        RECT 235.665 64.365 235.835 64.535 ;
        RECT 236.025 64.365 236.195 64.535 ;
        RECT 236.385 64.365 236.555 64.535 ;
        RECT 236.745 64.365 236.915 64.535 ;
        RECT 237.105 64.365 237.275 64.535 ;
        RECT 237.465 64.365 237.635 64.535 ;
        RECT 237.825 64.365 237.995 64.535 ;
        RECT 238.185 64.365 238.355 64.535 ;
        RECT 238.545 64.365 238.715 64.535 ;
        RECT 238.905 64.365 239.075 64.535 ;
        RECT 239.265 64.365 239.435 64.535 ;
        RECT 239.625 64.365 239.795 64.535 ;
        RECT 239.985 64.365 240.155 64.535 ;
        RECT 240.345 64.365 240.515 64.535 ;
        RECT 240.705 64.365 240.875 64.535 ;
        RECT 241.065 64.365 241.235 64.535 ;
        RECT 241.425 64.365 241.595 64.535 ;
        RECT 241.785 64.365 241.955 64.535 ;
        RECT 242.145 64.365 242.315 64.535 ;
        RECT 242.505 64.365 242.675 64.535 ;
        RECT 242.865 64.365 243.035 64.535 ;
        RECT 243.225 64.365 243.395 64.535 ;
        RECT 243.585 64.365 243.755 64.535 ;
        RECT 243.945 64.365 244.115 64.535 ;
        RECT 244.305 64.365 244.475 64.535 ;
        RECT 244.665 64.365 244.835 64.535 ;
        RECT 245.025 64.365 245.195 64.535 ;
        RECT 245.385 64.365 245.555 64.535 ;
        RECT 245.745 64.365 245.915 64.535 ;
        RECT 246.105 64.365 246.275 64.535 ;
        RECT 246.465 64.365 246.635 64.535 ;
        RECT 246.825 64.365 246.995 64.535 ;
        RECT 247.185 64.365 247.355 64.535 ;
        RECT 247.545 64.365 247.715 64.535 ;
        RECT 247.905 64.365 248.075 64.535 ;
        RECT 248.265 64.365 248.435 64.535 ;
        RECT 248.625 64.365 248.795 64.535 ;
        RECT 248.985 64.365 249.155 64.535 ;
        RECT 249.345 64.365 249.515 64.535 ;
        RECT 249.705 64.365 249.875 64.535 ;
        RECT 250.065 64.365 250.235 64.535 ;
        RECT 250.425 64.365 250.595 64.535 ;
        RECT 251.540 64.375 251.710 64.545 ;
        RECT 251.900 64.375 252.070 64.545 ;
        RECT 252.260 64.375 252.430 64.545 ;
        RECT 252.620 64.375 252.790 64.545 ;
        RECT 252.980 64.375 253.150 64.545 ;
        RECT 253.340 64.375 253.510 64.545 ;
        RECT 253.700 64.375 253.870 64.545 ;
        RECT 254.060 64.375 254.230 64.545 ;
        RECT 254.420 64.375 254.590 64.545 ;
        RECT 254.780 64.375 254.950 64.545 ;
        RECT 255.140 64.375 255.310 64.545 ;
        RECT 255.500 64.375 255.670 64.545 ;
        RECT 255.860 64.375 256.030 64.545 ;
        RECT 334.680 64.925 334.850 65.095 ;
        RECT 282.105 64.425 282.275 64.595 ;
        RECT 282.465 64.425 282.635 64.595 ;
        RECT 282.825 64.425 282.995 64.595 ;
        RECT 283.185 64.425 283.355 64.595 ;
        RECT 283.545 64.425 283.715 64.595 ;
        RECT 283.905 64.425 284.075 64.595 ;
        RECT 284.265 64.425 284.435 64.595 ;
        RECT 284.625 64.425 284.795 64.595 ;
        RECT 284.985 64.425 285.155 64.595 ;
        RECT 285.345 64.425 285.515 64.595 ;
        RECT 285.705 64.425 285.875 64.595 ;
        RECT 286.065 64.425 286.235 64.595 ;
        RECT 286.425 64.425 286.595 64.595 ;
        RECT 286.785 64.425 286.955 64.595 ;
        RECT 287.145 64.425 287.315 64.595 ;
        RECT 287.505 64.425 287.675 64.595 ;
        RECT 287.865 64.425 288.035 64.595 ;
        RECT 288.225 64.425 288.395 64.595 ;
        RECT 288.585 64.425 288.755 64.595 ;
        RECT 288.945 64.425 289.115 64.595 ;
        RECT 289.305 64.425 289.475 64.595 ;
        RECT 289.665 64.425 289.835 64.595 ;
        RECT 290.025 64.425 290.195 64.595 ;
        RECT 290.385 64.425 290.555 64.595 ;
        RECT 290.745 64.425 290.915 64.595 ;
        RECT 291.105 64.425 291.275 64.595 ;
        RECT 291.465 64.425 291.635 64.595 ;
        RECT 291.825 64.425 291.995 64.595 ;
        RECT 292.185 64.425 292.355 64.595 ;
        RECT 292.545 64.425 292.715 64.595 ;
        RECT 292.905 64.425 293.075 64.595 ;
        RECT 293.265 64.425 293.435 64.595 ;
        RECT 293.625 64.425 293.795 64.595 ;
        RECT 293.985 64.425 294.155 64.595 ;
        RECT 294.345 64.425 294.515 64.595 ;
        RECT 294.705 64.425 294.875 64.595 ;
        RECT 295.065 64.425 295.235 64.595 ;
        RECT 295.425 64.425 295.595 64.595 ;
        RECT 295.785 64.425 295.955 64.595 ;
        RECT 296.145 64.425 296.315 64.595 ;
        RECT 296.505 64.425 296.675 64.595 ;
        RECT 296.865 64.425 297.035 64.595 ;
        RECT 297.225 64.425 297.395 64.595 ;
        RECT 297.585 64.425 297.755 64.595 ;
        RECT 297.945 64.425 298.115 64.595 ;
        RECT 298.305 64.425 298.475 64.595 ;
        RECT 298.665 64.425 298.835 64.595 ;
        RECT 299.025 64.425 299.195 64.595 ;
        RECT 299.385 64.425 299.555 64.595 ;
        RECT 299.745 64.425 299.915 64.595 ;
        RECT 300.105 64.425 300.275 64.595 ;
        RECT 300.465 64.425 300.635 64.595 ;
        RECT 300.825 64.425 300.995 64.595 ;
        RECT 301.185 64.425 301.355 64.595 ;
        RECT 301.545 64.425 301.715 64.595 ;
        RECT 301.905 64.425 302.075 64.595 ;
        RECT 302.265 64.425 302.435 64.595 ;
        RECT 302.625 64.425 302.795 64.595 ;
        RECT 302.985 64.425 303.155 64.595 ;
        RECT 303.345 64.425 303.515 64.595 ;
        RECT 303.705 64.425 303.875 64.595 ;
        RECT 304.065 64.425 304.235 64.595 ;
        RECT 304.425 64.425 304.595 64.595 ;
        RECT 304.785 64.425 304.955 64.595 ;
        RECT 305.145 64.425 305.315 64.595 ;
        RECT 305.505 64.425 305.675 64.595 ;
        RECT 305.865 64.425 306.035 64.595 ;
        RECT 306.225 64.425 306.395 64.595 ;
        RECT 308.265 64.365 308.435 64.535 ;
        RECT 308.625 64.365 308.795 64.535 ;
        RECT 308.985 64.365 309.155 64.535 ;
        RECT 309.345 64.365 309.515 64.535 ;
        RECT 309.705 64.365 309.875 64.535 ;
        RECT 310.065 64.365 310.235 64.535 ;
        RECT 310.425 64.365 310.595 64.535 ;
        RECT 310.785 64.365 310.955 64.535 ;
        RECT 311.145 64.365 311.315 64.535 ;
        RECT 311.505 64.365 311.675 64.535 ;
        RECT 311.865 64.365 312.035 64.535 ;
        RECT 312.225 64.365 312.395 64.535 ;
        RECT 312.585 64.365 312.755 64.535 ;
        RECT 312.945 64.365 313.115 64.535 ;
        RECT 313.305 64.365 313.475 64.535 ;
        RECT 313.665 64.365 313.835 64.535 ;
        RECT 314.025 64.365 314.195 64.535 ;
        RECT 314.385 64.365 314.555 64.535 ;
        RECT 314.745 64.365 314.915 64.535 ;
        RECT 315.105 64.365 315.275 64.535 ;
        RECT 315.465 64.365 315.635 64.535 ;
        RECT 315.825 64.365 315.995 64.535 ;
        RECT 316.185 64.365 316.355 64.535 ;
        RECT 316.545 64.365 316.715 64.535 ;
        RECT 316.905 64.365 317.075 64.535 ;
        RECT 317.265 64.365 317.435 64.535 ;
        RECT 317.625 64.365 317.795 64.535 ;
        RECT 317.985 64.365 318.155 64.535 ;
        RECT 318.345 64.365 318.515 64.535 ;
        RECT 318.705 64.365 318.875 64.535 ;
        RECT 319.065 64.365 319.235 64.535 ;
        RECT 319.425 64.365 319.595 64.535 ;
        RECT 319.785 64.365 319.955 64.535 ;
        RECT 320.145 64.365 320.315 64.535 ;
        RECT 320.505 64.365 320.675 64.535 ;
        RECT 320.865 64.365 321.035 64.535 ;
        RECT 321.225 64.365 321.395 64.535 ;
        RECT 321.585 64.365 321.755 64.535 ;
        RECT 321.945 64.365 322.115 64.535 ;
        RECT 322.305 64.365 322.475 64.535 ;
        RECT 322.665 64.365 322.835 64.535 ;
        RECT 323.025 64.365 323.195 64.535 ;
        RECT 323.385 64.365 323.555 64.535 ;
        RECT 323.745 64.365 323.915 64.535 ;
        RECT 324.105 64.365 324.275 64.535 ;
        RECT 324.465 64.365 324.635 64.535 ;
        RECT 324.825 64.365 324.995 64.535 ;
        RECT 325.185 64.365 325.355 64.535 ;
        RECT 325.545 64.365 325.715 64.535 ;
        RECT 325.905 64.365 326.075 64.535 ;
        RECT 326.265 64.365 326.435 64.535 ;
        RECT 326.625 64.365 326.795 64.535 ;
        RECT 326.985 64.365 327.155 64.535 ;
        RECT 327.345 64.365 327.515 64.535 ;
        RECT 327.705 64.365 327.875 64.535 ;
      LAYER met1 ;
        RECT 209.230 133.210 278.240 134.030 ;
        RECT 308.095 133.800 328.000 133.815 ;
        RECT 308.095 133.795 332.435 133.800 ;
        RECT 308.035 133.365 332.435 133.795 ;
        RECT 308.035 133.360 328.060 133.365 ;
        RECT 308.095 133.340 328.000 133.360 ;
        RECT 202.580 65.070 203.315 131.540 ;
        RECT 330.225 131.200 332.385 133.365 ;
        RECT 264.275 96.635 264.740 99.285 ;
        RECT 264.220 96.065 265.400 96.245 ;
        RECT 264.220 95.955 265.495 96.065 ;
        RECT 263.155 95.725 265.495 95.955 ;
        RECT 263.155 95.590 263.575 95.725 ;
        RECT 264.220 95.630 265.495 95.725 ;
        RECT 264.220 95.330 265.400 95.630 ;
        RECT 264.245 92.860 265.425 93.090 ;
        RECT 264.235 92.750 265.490 92.860 ;
        RECT 263.160 92.740 265.490 92.750 ;
        RECT 263.155 92.520 265.490 92.740 ;
        RECT 263.155 92.510 263.575 92.520 ;
        RECT 264.235 92.425 265.490 92.520 ;
        RECT 264.245 92.175 265.425 92.425 ;
        RECT 264.285 89.855 265.465 90.075 ;
        RECT 264.240 89.765 265.495 89.855 ;
        RECT 263.170 89.660 265.495 89.765 ;
        RECT 263.155 89.535 265.495 89.660 ;
        RECT 263.155 89.430 263.575 89.535 ;
        RECT 264.240 89.420 265.495 89.535 ;
        RECT 264.285 89.160 265.465 89.420 ;
        RECT 258.465 84.230 258.935 85.820 ;
        RECT 263.155 85.605 263.575 85.790 ;
        RECT 264.275 85.715 265.455 85.955 ;
        RECT 264.250 85.605 265.505 85.715 ;
        RECT 266.185 85.605 266.605 85.790 ;
        RECT 263.155 85.560 266.640 85.605 ;
        RECT 263.175 85.360 266.640 85.560 ;
        RECT 264.250 85.280 265.505 85.360 ;
        RECT 264.275 85.040 265.455 85.280 ;
        RECT 267.140 79.740 270.900 80.370 ;
        RECT 266.555 78.480 266.975 78.510 ;
        RECT 266.550 78.220 266.980 78.480 ;
        RECT 267.885 78.220 270.155 79.740 ;
        RECT 271.065 78.480 271.485 78.510 ;
        RECT 271.060 78.220 271.490 78.480 ;
        RECT 266.550 76.330 271.490 78.220 ;
        RECT 266.550 76.010 266.980 76.330 ;
        RECT 266.555 75.990 266.975 76.010 ;
        RECT 267.885 74.740 270.155 76.330 ;
        RECT 271.060 76.010 271.490 76.330 ;
        RECT 271.065 75.990 271.485 76.010 ;
        RECT 267.290 74.110 270.750 74.740 ;
        RECT 267.365 73.520 270.745 74.110 ;
        RECT 255.835 73.515 281.445 73.520 ;
        RECT 255.835 72.395 281.495 73.515 ;
        RECT 205.385 65.070 207.545 66.910 ;
        RECT 255.835 65.070 256.940 72.395 ;
        RECT 202.575 63.965 256.940 65.070 ;
        RECT 280.740 64.835 281.495 72.395 ;
        RECT 334.200 64.835 335.215 133.975 ;
        RECT 280.740 64.080 335.215 64.835 ;
      LAYER via ;
        RECT 230.875 133.455 231.135 133.715 ;
        RECT 231.195 133.455 231.455 133.715 ;
        RECT 231.515 133.455 231.775 133.715 ;
        RECT 231.835 133.455 232.095 133.715 ;
        RECT 232.155 133.455 232.415 133.715 ;
        RECT 232.475 133.455 232.735 133.715 ;
        RECT 232.795 133.455 233.055 133.715 ;
        RECT 233.115 133.455 233.375 133.715 ;
        RECT 233.435 133.455 233.695 133.715 ;
        RECT 233.755 133.455 234.015 133.715 ;
        RECT 234.075 133.455 234.335 133.715 ;
        RECT 234.395 133.455 234.655 133.715 ;
        RECT 234.715 133.455 234.975 133.715 ;
        RECT 235.035 133.455 235.295 133.715 ;
        RECT 235.355 133.455 235.615 133.715 ;
        RECT 235.675 133.455 235.935 133.715 ;
        RECT 235.995 133.455 236.255 133.715 ;
        RECT 236.315 133.455 236.575 133.715 ;
        RECT 236.635 133.455 236.895 133.715 ;
        RECT 236.955 133.455 237.215 133.715 ;
        RECT 237.275 133.455 237.535 133.715 ;
        RECT 237.595 133.455 237.855 133.715 ;
        RECT 237.915 133.455 238.175 133.715 ;
        RECT 238.235 133.455 238.495 133.715 ;
        RECT 238.555 133.455 238.815 133.715 ;
        RECT 238.875 133.455 239.135 133.715 ;
        RECT 239.195 133.455 239.455 133.715 ;
        RECT 239.515 133.455 239.775 133.715 ;
        RECT 239.835 133.455 240.095 133.715 ;
        RECT 240.155 133.455 240.415 133.715 ;
        RECT 240.475 133.455 240.735 133.715 ;
        RECT 240.795 133.455 241.055 133.715 ;
        RECT 241.115 133.455 241.375 133.715 ;
        RECT 241.435 133.455 241.695 133.715 ;
        RECT 241.755 133.455 242.015 133.715 ;
        RECT 242.075 133.455 242.335 133.715 ;
        RECT 242.395 133.455 242.655 133.715 ;
        RECT 242.715 133.455 242.975 133.715 ;
        RECT 243.035 133.455 243.295 133.715 ;
        RECT 243.355 133.455 243.615 133.715 ;
        RECT 243.675 133.455 243.935 133.715 ;
        RECT 243.995 133.455 244.255 133.715 ;
        RECT 244.315 133.455 244.575 133.715 ;
        RECT 244.635 133.455 244.895 133.715 ;
        RECT 244.955 133.455 245.215 133.715 ;
        RECT 245.275 133.455 245.535 133.715 ;
        RECT 245.595 133.455 245.855 133.715 ;
        RECT 245.915 133.455 246.175 133.715 ;
        RECT 246.235 133.455 246.495 133.715 ;
        RECT 246.555 133.455 246.815 133.715 ;
        RECT 246.875 133.455 247.135 133.715 ;
        RECT 247.195 133.455 247.455 133.715 ;
        RECT 247.515 133.455 247.775 133.715 ;
        RECT 247.835 133.455 248.095 133.715 ;
        RECT 248.155 133.455 248.415 133.715 ;
        RECT 248.475 133.455 248.735 133.715 ;
        RECT 248.795 133.455 249.055 133.715 ;
        RECT 249.115 133.455 249.375 133.715 ;
        RECT 249.435 133.455 249.695 133.715 ;
        RECT 249.755 133.455 250.015 133.715 ;
        RECT 250.075 133.455 250.335 133.715 ;
        RECT 250.395 133.455 250.655 133.715 ;
        RECT 308.160 133.450 308.420 133.710 ;
        RECT 308.480 133.450 308.740 133.710 ;
        RECT 308.800 133.450 309.060 133.710 ;
        RECT 309.120 133.450 309.380 133.710 ;
        RECT 309.440 133.450 309.700 133.710 ;
        RECT 309.760 133.450 310.020 133.710 ;
        RECT 310.080 133.450 310.340 133.710 ;
        RECT 310.400 133.450 310.660 133.710 ;
        RECT 310.720 133.450 310.980 133.710 ;
        RECT 311.040 133.450 311.300 133.710 ;
        RECT 311.360 133.450 311.620 133.710 ;
        RECT 311.680 133.450 311.940 133.710 ;
        RECT 312.000 133.450 312.260 133.710 ;
        RECT 312.320 133.450 312.580 133.710 ;
        RECT 312.640 133.450 312.900 133.710 ;
        RECT 312.960 133.450 313.220 133.710 ;
        RECT 313.280 133.450 313.540 133.710 ;
        RECT 313.600 133.450 313.860 133.710 ;
        RECT 313.920 133.450 314.180 133.710 ;
        RECT 314.240 133.450 314.500 133.710 ;
        RECT 314.560 133.450 314.820 133.710 ;
        RECT 314.880 133.450 315.140 133.710 ;
        RECT 315.200 133.450 315.460 133.710 ;
        RECT 315.520 133.450 315.780 133.710 ;
        RECT 315.840 133.450 316.100 133.710 ;
        RECT 316.160 133.450 316.420 133.710 ;
        RECT 316.480 133.450 316.740 133.710 ;
        RECT 316.800 133.450 317.060 133.710 ;
        RECT 317.120 133.450 317.380 133.710 ;
        RECT 317.440 133.450 317.700 133.710 ;
        RECT 317.760 133.450 318.020 133.710 ;
        RECT 318.080 133.450 318.340 133.710 ;
        RECT 318.400 133.450 318.660 133.710 ;
        RECT 318.720 133.450 318.980 133.710 ;
        RECT 319.040 133.450 319.300 133.710 ;
        RECT 319.360 133.450 319.620 133.710 ;
        RECT 319.680 133.450 319.940 133.710 ;
        RECT 320.000 133.450 320.260 133.710 ;
        RECT 320.320 133.450 320.580 133.710 ;
        RECT 320.640 133.450 320.900 133.710 ;
        RECT 320.960 133.450 321.220 133.710 ;
        RECT 321.280 133.450 321.540 133.710 ;
        RECT 321.600 133.450 321.860 133.710 ;
        RECT 321.920 133.450 322.180 133.710 ;
        RECT 322.240 133.450 322.500 133.710 ;
        RECT 322.560 133.450 322.820 133.710 ;
        RECT 322.880 133.450 323.140 133.710 ;
        RECT 323.200 133.450 323.460 133.710 ;
        RECT 323.520 133.450 323.780 133.710 ;
        RECT 323.840 133.450 324.100 133.710 ;
        RECT 324.160 133.450 324.420 133.710 ;
        RECT 324.480 133.450 324.740 133.710 ;
        RECT 324.800 133.450 325.060 133.710 ;
        RECT 325.120 133.450 325.380 133.710 ;
        RECT 325.440 133.450 325.700 133.710 ;
        RECT 325.760 133.450 326.020 133.710 ;
        RECT 326.080 133.450 326.340 133.710 ;
        RECT 326.400 133.450 326.660 133.710 ;
        RECT 326.720 133.450 326.980 133.710 ;
        RECT 327.040 133.450 327.300 133.710 ;
        RECT 327.360 133.450 327.620 133.710 ;
        RECT 327.680 133.450 327.940 133.710 ;
        RECT 264.380 98.950 264.640 99.210 ;
        RECT 264.380 98.630 264.640 98.890 ;
        RECT 264.380 98.310 264.640 98.570 ;
        RECT 264.380 97.990 264.640 98.250 ;
        RECT 264.380 97.670 264.640 97.930 ;
        RECT 264.380 97.350 264.640 97.610 ;
        RECT 264.380 97.030 264.640 97.290 ;
        RECT 264.380 96.710 264.640 96.970 ;
        RECT 264.360 95.500 265.260 96.080 ;
        RECT 264.385 92.345 265.285 92.925 ;
        RECT 264.425 89.330 265.325 89.910 ;
        RECT 258.570 85.495 258.830 85.755 ;
        RECT 258.570 85.175 258.830 85.435 ;
        RECT 258.570 84.855 258.830 85.115 ;
        RECT 264.415 85.210 265.315 85.790 ;
        RECT 258.570 84.535 258.830 84.795 ;
        RECT 230.900 64.320 231.160 64.580 ;
        RECT 231.220 64.320 231.480 64.580 ;
        RECT 231.540 64.320 231.800 64.580 ;
        RECT 231.860 64.320 232.120 64.580 ;
        RECT 232.180 64.320 232.440 64.580 ;
        RECT 232.500 64.320 232.760 64.580 ;
        RECT 232.820 64.320 233.080 64.580 ;
        RECT 233.140 64.320 233.400 64.580 ;
        RECT 233.460 64.320 233.720 64.580 ;
        RECT 233.780 64.320 234.040 64.580 ;
        RECT 234.100 64.320 234.360 64.580 ;
        RECT 234.420 64.320 234.680 64.580 ;
        RECT 234.740 64.320 235.000 64.580 ;
        RECT 235.060 64.320 235.320 64.580 ;
        RECT 235.380 64.320 235.640 64.580 ;
        RECT 235.700 64.320 235.960 64.580 ;
        RECT 236.020 64.320 236.280 64.580 ;
        RECT 236.340 64.320 236.600 64.580 ;
        RECT 236.660 64.320 236.920 64.580 ;
        RECT 236.980 64.320 237.240 64.580 ;
        RECT 237.300 64.320 237.560 64.580 ;
        RECT 237.620 64.320 237.880 64.580 ;
        RECT 237.940 64.320 238.200 64.580 ;
        RECT 238.260 64.320 238.520 64.580 ;
        RECT 238.580 64.320 238.840 64.580 ;
        RECT 238.900 64.320 239.160 64.580 ;
        RECT 239.220 64.320 239.480 64.580 ;
        RECT 239.540 64.320 239.800 64.580 ;
        RECT 239.860 64.320 240.120 64.580 ;
        RECT 240.180 64.320 240.440 64.580 ;
        RECT 240.500 64.320 240.760 64.580 ;
        RECT 240.820 64.320 241.080 64.580 ;
        RECT 241.140 64.320 241.400 64.580 ;
        RECT 241.460 64.320 241.720 64.580 ;
        RECT 241.780 64.320 242.040 64.580 ;
        RECT 242.100 64.320 242.360 64.580 ;
        RECT 242.420 64.320 242.680 64.580 ;
        RECT 242.740 64.320 243.000 64.580 ;
        RECT 243.060 64.320 243.320 64.580 ;
        RECT 243.380 64.320 243.640 64.580 ;
        RECT 243.700 64.320 243.960 64.580 ;
        RECT 244.020 64.320 244.280 64.580 ;
        RECT 244.340 64.320 244.600 64.580 ;
        RECT 244.660 64.320 244.920 64.580 ;
        RECT 244.980 64.320 245.240 64.580 ;
        RECT 245.300 64.320 245.560 64.580 ;
        RECT 245.620 64.320 245.880 64.580 ;
        RECT 245.940 64.320 246.200 64.580 ;
        RECT 246.260 64.320 246.520 64.580 ;
        RECT 246.580 64.320 246.840 64.580 ;
        RECT 246.900 64.320 247.160 64.580 ;
        RECT 247.220 64.320 247.480 64.580 ;
        RECT 247.540 64.320 247.800 64.580 ;
        RECT 247.860 64.320 248.120 64.580 ;
        RECT 248.180 64.320 248.440 64.580 ;
        RECT 248.500 64.320 248.760 64.580 ;
        RECT 248.820 64.320 249.080 64.580 ;
        RECT 249.140 64.320 249.400 64.580 ;
        RECT 249.460 64.320 249.720 64.580 ;
        RECT 249.780 64.320 250.040 64.580 ;
        RECT 250.100 64.320 250.360 64.580 ;
        RECT 250.420 64.320 250.680 64.580 ;
        RECT 308.180 64.320 308.440 64.580 ;
        RECT 308.500 64.320 308.760 64.580 ;
        RECT 308.820 64.320 309.080 64.580 ;
        RECT 309.140 64.320 309.400 64.580 ;
        RECT 309.460 64.320 309.720 64.580 ;
        RECT 309.780 64.320 310.040 64.580 ;
        RECT 310.100 64.320 310.360 64.580 ;
        RECT 310.420 64.320 310.680 64.580 ;
        RECT 310.740 64.320 311.000 64.580 ;
        RECT 311.060 64.320 311.320 64.580 ;
        RECT 311.380 64.320 311.640 64.580 ;
        RECT 311.700 64.320 311.960 64.580 ;
        RECT 312.020 64.320 312.280 64.580 ;
        RECT 312.340 64.320 312.600 64.580 ;
        RECT 312.660 64.320 312.920 64.580 ;
        RECT 312.980 64.320 313.240 64.580 ;
        RECT 313.300 64.320 313.560 64.580 ;
        RECT 313.620 64.320 313.880 64.580 ;
        RECT 313.940 64.320 314.200 64.580 ;
        RECT 314.260 64.320 314.520 64.580 ;
        RECT 314.580 64.320 314.840 64.580 ;
        RECT 314.900 64.320 315.160 64.580 ;
        RECT 315.220 64.320 315.480 64.580 ;
        RECT 315.540 64.320 315.800 64.580 ;
        RECT 315.860 64.320 316.120 64.580 ;
        RECT 316.180 64.320 316.440 64.580 ;
        RECT 316.500 64.320 316.760 64.580 ;
        RECT 316.820 64.320 317.080 64.580 ;
        RECT 317.140 64.320 317.400 64.580 ;
        RECT 317.460 64.320 317.720 64.580 ;
        RECT 317.780 64.320 318.040 64.580 ;
        RECT 318.100 64.320 318.360 64.580 ;
        RECT 318.420 64.320 318.680 64.580 ;
        RECT 318.740 64.320 319.000 64.580 ;
        RECT 319.060 64.320 319.320 64.580 ;
        RECT 319.380 64.320 319.640 64.580 ;
        RECT 319.700 64.320 319.960 64.580 ;
        RECT 320.020 64.320 320.280 64.580 ;
        RECT 320.340 64.320 320.600 64.580 ;
        RECT 320.660 64.320 320.920 64.580 ;
        RECT 320.980 64.320 321.240 64.580 ;
        RECT 321.300 64.320 321.560 64.580 ;
        RECT 321.620 64.320 321.880 64.580 ;
        RECT 321.940 64.320 322.200 64.580 ;
        RECT 322.260 64.320 322.520 64.580 ;
        RECT 322.580 64.320 322.840 64.580 ;
        RECT 322.900 64.320 323.160 64.580 ;
        RECT 323.220 64.320 323.480 64.580 ;
        RECT 323.540 64.320 323.800 64.580 ;
        RECT 323.860 64.320 324.120 64.580 ;
        RECT 324.180 64.320 324.440 64.580 ;
        RECT 324.500 64.320 324.760 64.580 ;
        RECT 324.820 64.320 325.080 64.580 ;
        RECT 325.140 64.320 325.400 64.580 ;
        RECT 325.460 64.320 325.720 64.580 ;
        RECT 325.780 64.320 326.040 64.580 ;
        RECT 326.100 64.320 326.360 64.580 ;
        RECT 326.420 64.320 326.680 64.580 ;
        RECT 326.740 64.320 327.000 64.580 ;
        RECT 327.060 64.320 327.320 64.580 ;
        RECT 327.380 64.320 327.640 64.580 ;
        RECT 327.700 64.320 327.960 64.580 ;
      LAYER met2 ;
        RECT 230.755 100.810 250.755 134.100 ;
        RECT 308.055 133.765 328.055 134.100 ;
        RECT 308.045 133.390 328.055 133.765 ;
        RECT 230.755 94.780 265.910 100.810 ;
        RECT 230.755 89.925 250.755 94.780 ;
        RECT 263.675 89.925 265.910 94.780 ;
        RECT 230.755 84.530 265.910 89.925 ;
        RECT 230.755 83.895 256.720 84.530 ;
        RECT 230.755 63.930 250.755 83.895 ;
        RECT 308.055 63.930 328.055 133.390 ;
      LAYER via2 ;
        RECT 235.220 132.565 236.700 134.000 ;
        RECT 238.550 132.565 240.030 134.000 ;
        RECT 241.845 132.545 243.325 133.980 ;
        RECT 245.160 132.545 246.640 133.980 ;
        RECT 312.405 132.565 313.885 134.000 ;
        RECT 315.735 132.565 317.215 134.000 ;
        RECT 319.030 132.545 320.510 133.980 ;
        RECT 322.345 132.545 323.825 133.980 ;
        RECT 235.220 64.105 236.700 65.540 ;
        RECT 238.550 64.105 240.030 65.540 ;
        RECT 241.845 64.085 243.325 65.520 ;
        RECT 245.160 64.085 246.640 65.520 ;
        RECT 312.405 64.105 313.885 65.540 ;
        RECT 315.735 64.105 317.215 65.540 ;
        RECT 319.030 64.085 320.510 65.520 ;
        RECT 322.345 64.085 323.825 65.520 ;
      LAYER met3 ;
        RECT 230.755 132.390 250.755 134.100 ;
        RECT 307.940 132.390 327.940 134.100 ;
        RECT 230.755 63.930 250.755 65.640 ;
        RECT 307.940 63.930 327.940 65.640 ;
      LAYER via3 ;
        RECT 235.200 132.545 236.720 134.020 ;
        RECT 238.530 132.545 240.050 134.020 ;
        RECT 241.825 132.525 243.345 134.000 ;
        RECT 245.140 132.525 246.660 134.000 ;
        RECT 312.385 132.545 313.905 134.020 ;
        RECT 315.715 132.545 317.235 134.020 ;
        RECT 319.010 132.525 320.530 134.000 ;
        RECT 322.325 132.525 323.845 134.000 ;
        RECT 235.200 64.085 236.720 65.560 ;
        RECT 238.530 64.085 240.050 65.560 ;
        RECT 241.825 64.065 243.345 65.540 ;
        RECT 245.140 64.065 246.660 65.540 ;
        RECT 312.385 64.085 313.905 65.560 ;
        RECT 315.715 64.085 317.235 65.560 ;
        RECT 319.010 64.065 320.530 65.540 ;
        RECT 322.325 64.065 323.845 65.540 ;
      LAYER met4 ;
        RECT 235.165 3.300 236.765 211.800 ;
        RECT 238.465 3.300 240.065 211.800 ;
        RECT 241.765 3.300 243.365 211.800 ;
        RECT 245.065 3.300 246.665 211.800 ;
        RECT 312.350 3.300 313.950 211.800 ;
        RECT 315.650 3.300 317.250 211.800 ;
        RECT 318.950 3.300 320.550 211.800 ;
        RECT 322.250 3.300 323.850 211.800 ;
    END
  END vdda1
  PIN vssa1
    ANTENNADIFFAREA 167.107590 ;
    PORT
      LAYER pwell ;
        RECT 204.555 131.680 255.275 132.110 ;
        RECT 204.555 84.150 204.985 131.680 ;
        RECT 254.845 84.150 255.275 131.680 ;
        RECT 282.445 131.900 333.165 132.330 ;
        RECT 256.615 131.100 281.335 131.530 ;
        RECT 256.615 102.800 257.045 131.100 ;
        RECT 280.905 102.800 281.335 131.100 ;
        RECT 256.615 102.370 281.335 102.800 ;
        RECT 269.235 97.530 271.825 100.210 ;
        RECT 272.235 97.530 274.825 100.210 ;
        RECT 269.235 94.750 271.825 97.430 ;
        RECT 272.235 94.750 274.825 97.430 ;
        RECT 269.235 91.970 271.825 94.650 ;
        RECT 272.235 91.970 274.825 94.650 ;
        RECT 275.865 91.960 278.455 94.640 ;
        RECT 269.235 89.190 271.825 91.870 ;
        RECT 272.235 89.190 274.825 91.870 ;
        RECT 275.865 89.180 278.455 91.860 ;
        RECT 257.080 87.435 258.810 89.165 ;
        RECT 204.555 83.720 255.275 84.150 ;
        RECT 256.375 86.155 259.485 86.585 ;
        RECT 269.235 86.410 271.825 89.090 ;
        RECT 272.235 86.410 274.825 89.090 ;
        RECT 275.865 86.400 278.455 89.080 ;
        RECT 256.375 83.905 256.805 86.155 ;
        RECT 259.055 83.905 259.485 86.155 ;
        RECT 256.375 83.475 259.485 83.905 ;
        RECT 269.235 83.630 271.825 86.310 ;
        RECT 272.235 83.630 274.825 86.310 ;
        RECT 275.865 83.620 278.455 86.300 ;
        RECT 204.605 82.200 255.325 82.630 ;
        RECT 204.605 66.210 205.035 82.200 ;
        RECT 254.895 66.210 255.325 82.200 ;
        RECT 258.470 77.440 261.370 80.120 ;
        RECT 276.670 77.440 279.570 80.120 ;
        RECT 258.460 74.410 261.360 77.090 ;
        RECT 276.680 74.410 279.580 77.090 ;
        RECT 204.605 65.780 255.325 66.210 ;
        RECT 282.445 66.110 282.875 131.900 ;
        RECT 332.735 66.110 333.165 131.900 ;
        RECT 282.445 65.680 333.165 66.110 ;
      LAYER li1 ;
        RECT 286.585 132.200 306.465 132.260 ;
        RECT 282.575 132.030 333.035 132.200 ;
        RECT 209.375 131.980 229.190 131.985 ;
        RECT 204.685 131.810 255.145 131.980 ;
        RECT 204.685 84.020 204.855 131.810 ;
        RECT 254.975 89.030 255.145 131.810 ;
        RECT 257.855 131.400 278.515 131.565 ;
        RECT 256.745 131.230 281.205 131.400 ;
        RECT 256.745 102.670 256.915 131.230 ;
        RECT 257.855 131.200 278.515 131.230 ;
        RECT 281.035 102.670 281.205 131.230 ;
        RECT 256.745 102.500 281.205 102.670 ;
        RECT 268.925 100.020 269.520 100.045 ;
        RECT 271.490 100.020 272.480 100.050 ;
        RECT 274.495 100.020 276.180 100.075 ;
        RECT 268.925 99.850 276.180 100.020 ;
        RECT 268.925 97.890 269.595 99.850 ;
        RECT 271.465 97.890 272.595 99.850 ;
        RECT 273.145 98.390 273.605 98.560 ;
        RECT 274.465 97.890 276.180 99.850 ;
        RECT 268.925 97.070 276.180 97.890 ;
        RECT 268.925 95.110 269.595 97.070 ;
        RECT 271.465 95.110 272.595 97.070 ;
        RECT 273.145 95.610 273.605 95.780 ;
        RECT 274.465 95.110 276.180 97.070 ;
        RECT 268.925 94.450 276.180 95.110 ;
        RECT 268.925 94.290 278.265 94.450 ;
        RECT 268.925 92.330 269.595 94.290 ;
        RECT 271.465 92.330 272.595 94.290 ;
        RECT 274.465 94.280 278.265 94.290 ;
        RECT 273.145 92.830 273.605 93.000 ;
        RECT 274.465 92.330 276.225 94.280 ;
        RECT 276.775 92.820 277.235 92.990 ;
        RECT 268.925 92.320 276.225 92.330 ;
        RECT 278.095 92.320 278.265 94.280 ;
        RECT 268.925 91.510 278.265 92.320 ;
        RECT 268.925 89.550 269.595 91.510 ;
        RECT 271.465 89.550 272.595 91.510 ;
        RECT 274.465 91.500 278.265 91.510 ;
        RECT 273.145 90.050 273.605 90.220 ;
        RECT 274.465 89.550 276.225 91.500 ;
        RECT 276.775 90.830 277.235 91.000 ;
        RECT 268.925 89.540 276.225 89.550 ;
        RECT 278.095 89.540 278.265 91.500 ;
        RECT 268.925 89.370 278.265 89.540 ;
        RECT 257.210 89.030 258.680 89.035 ;
        RECT 254.975 88.865 258.990 89.030 ;
        RECT 254.975 87.735 257.380 88.865 ;
        RECT 258.500 87.735 258.990 88.865 ;
        RECT 254.975 87.670 258.990 87.735 ;
        RECT 268.925 88.890 278.250 89.370 ;
        RECT 268.925 88.730 278.265 88.890 ;
        RECT 254.975 87.115 258.995 87.670 ;
        RECT 254.975 86.285 259.515 87.115 ;
        RECT 209.470 84.020 229.285 84.060 ;
        RECT 254.975 84.020 256.675 86.285 ;
        RECT 204.685 83.850 256.675 84.020 ;
        RECT 209.470 83.800 229.285 83.850 ;
        RECT 256.505 83.775 256.675 83.850 ;
        RECT 259.175 83.775 259.515 86.285 ;
        RECT 268.925 86.770 269.595 88.730 ;
        RECT 271.465 86.770 272.595 88.730 ;
        RECT 274.465 88.720 278.265 88.730 ;
        RECT 273.145 87.270 273.605 87.440 ;
        RECT 274.465 86.770 276.225 88.720 ;
        RECT 276.775 87.260 277.235 87.430 ;
        RECT 268.925 86.760 276.225 86.770 ;
        RECT 278.095 86.760 278.265 88.720 ;
        RECT 268.925 86.590 278.265 86.760 ;
        RECT 268.925 86.110 278.250 86.590 ;
        RECT 268.925 85.950 278.265 86.110 ;
        RECT 268.925 83.990 269.595 85.950 ;
        RECT 271.465 83.990 272.595 85.950 ;
        RECT 274.465 85.940 278.265 85.950 ;
        RECT 273.145 84.490 273.605 84.660 ;
        RECT 274.465 83.990 276.225 85.940 ;
        RECT 268.925 83.980 276.225 83.990 ;
        RECT 278.095 83.980 278.265 85.940 ;
        RECT 268.925 83.845 278.265 83.980 ;
        RECT 268.925 83.840 271.635 83.845 ;
        RECT 269.425 83.820 271.635 83.840 ;
        RECT 272.425 83.830 278.265 83.845 ;
        RECT 272.425 83.820 274.635 83.830 ;
        RECT 276.055 83.810 278.265 83.830 ;
        RECT 256.505 83.605 259.515 83.775 ;
        RECT 209.470 82.500 229.285 82.545 ;
        RECT 204.735 82.330 255.195 82.500 ;
        RECT 204.735 66.080 204.905 82.330 ;
        RECT 209.470 82.285 229.285 82.330 ;
        RECT 209.445 66.080 229.260 66.120 ;
        RECT 255.025 66.080 255.195 82.330 ;
        RECT 258.020 79.740 261.510 80.370 ;
        RECT 258.020 77.810 258.850 79.740 ;
        RECT 259.690 79.090 260.150 79.260 ;
        RECT 260.980 77.810 261.510 79.740 ;
        RECT 258.020 76.730 261.510 77.810 ;
        RECT 258.020 74.790 258.850 76.730 ;
        RECT 259.680 75.270 260.140 75.440 ;
        RECT 260.980 74.790 261.510 76.730 ;
        RECT 258.020 74.160 261.510 74.790 ;
        RECT 276.530 79.740 280.020 80.370 ;
        RECT 276.530 77.810 277.060 79.740 ;
        RECT 277.890 79.090 278.350 79.260 ;
        RECT 279.190 77.810 280.020 79.740 ;
        RECT 276.530 76.730 280.020 77.810 ;
        RECT 276.530 74.790 277.060 76.730 ;
        RECT 277.900 75.270 278.360 75.440 ;
        RECT 279.190 74.790 280.020 76.730 ;
        RECT 276.530 74.160 280.020 74.790 ;
        RECT 204.735 65.910 255.195 66.080 ;
        RECT 282.575 65.980 282.745 132.030 ;
        RECT 286.585 132.000 306.465 132.030 ;
        RECT 286.595 65.980 306.475 66.030 ;
        RECT 332.865 65.980 333.035 132.030 ;
        RECT 209.445 65.860 229.260 65.910 ;
        RECT 282.575 65.810 333.035 65.980 ;
        RECT 286.595 65.770 306.475 65.810 ;
      LAYER mcon ;
        RECT 286.720 132.045 286.890 132.215 ;
        RECT 287.080 132.045 287.250 132.215 ;
        RECT 287.440 132.045 287.610 132.215 ;
        RECT 287.800 132.045 287.970 132.215 ;
        RECT 288.160 132.045 288.330 132.215 ;
        RECT 288.520 132.045 288.690 132.215 ;
        RECT 288.880 132.045 289.050 132.215 ;
        RECT 289.240 132.045 289.410 132.215 ;
        RECT 289.600 132.045 289.770 132.215 ;
        RECT 289.960 132.045 290.130 132.215 ;
        RECT 290.320 132.045 290.490 132.215 ;
        RECT 290.680 132.045 290.850 132.215 ;
        RECT 291.040 132.045 291.210 132.215 ;
        RECT 291.400 132.045 291.570 132.215 ;
        RECT 291.760 132.045 291.930 132.215 ;
        RECT 292.120 132.045 292.290 132.215 ;
        RECT 292.480 132.045 292.650 132.215 ;
        RECT 292.840 132.045 293.010 132.215 ;
        RECT 293.200 132.045 293.370 132.215 ;
        RECT 293.560 132.045 293.730 132.215 ;
        RECT 293.920 132.045 294.090 132.215 ;
        RECT 294.280 132.045 294.450 132.215 ;
        RECT 294.640 132.045 294.810 132.215 ;
        RECT 295.000 132.045 295.170 132.215 ;
        RECT 295.360 132.045 295.530 132.215 ;
        RECT 295.720 132.045 295.890 132.215 ;
        RECT 296.080 132.045 296.250 132.215 ;
        RECT 296.440 132.045 296.610 132.215 ;
        RECT 296.800 132.045 296.970 132.215 ;
        RECT 297.160 132.045 297.330 132.215 ;
        RECT 297.520 132.045 297.690 132.215 ;
        RECT 297.880 132.045 298.050 132.215 ;
        RECT 298.240 132.045 298.410 132.215 ;
        RECT 298.600 132.045 298.770 132.215 ;
        RECT 298.960 132.045 299.130 132.215 ;
        RECT 299.320 132.045 299.490 132.215 ;
        RECT 299.680 132.045 299.850 132.215 ;
        RECT 300.040 132.045 300.210 132.215 ;
        RECT 300.400 132.045 300.570 132.215 ;
        RECT 300.760 132.045 300.930 132.215 ;
        RECT 301.120 132.045 301.290 132.215 ;
        RECT 301.480 132.045 301.650 132.215 ;
        RECT 301.840 132.045 302.010 132.215 ;
        RECT 302.200 132.045 302.370 132.215 ;
        RECT 302.560 132.045 302.730 132.215 ;
        RECT 302.920 132.045 303.090 132.215 ;
        RECT 303.280 132.045 303.450 132.215 ;
        RECT 303.640 132.045 303.810 132.215 ;
        RECT 304.000 132.045 304.170 132.215 ;
        RECT 304.360 132.045 304.530 132.215 ;
        RECT 304.720 132.045 304.890 132.215 ;
        RECT 305.080 132.045 305.250 132.215 ;
        RECT 305.440 132.045 305.610 132.215 ;
        RECT 305.800 132.045 305.970 132.215 ;
        RECT 306.160 132.045 306.330 132.215 ;
        RECT 209.480 131.815 209.650 131.985 ;
        RECT 209.840 131.815 210.010 131.985 ;
        RECT 210.200 131.815 210.370 131.985 ;
        RECT 210.560 131.815 210.730 131.985 ;
        RECT 210.920 131.815 211.090 131.985 ;
        RECT 211.280 131.815 211.450 131.985 ;
        RECT 211.640 131.815 211.810 131.985 ;
        RECT 212.000 131.815 212.170 131.985 ;
        RECT 212.360 131.815 212.530 131.985 ;
        RECT 212.720 131.815 212.890 131.985 ;
        RECT 213.080 131.815 213.250 131.985 ;
        RECT 213.440 131.815 213.610 131.985 ;
        RECT 213.800 131.815 213.970 131.985 ;
        RECT 214.160 131.815 214.330 131.985 ;
        RECT 214.520 131.815 214.690 131.985 ;
        RECT 214.880 131.815 215.050 131.985 ;
        RECT 215.240 131.815 215.410 131.985 ;
        RECT 215.600 131.815 215.770 131.985 ;
        RECT 215.960 131.815 216.130 131.985 ;
        RECT 216.320 131.815 216.490 131.985 ;
        RECT 216.680 131.815 216.850 131.985 ;
        RECT 217.040 131.815 217.210 131.985 ;
        RECT 217.400 131.815 217.570 131.985 ;
        RECT 217.760 131.815 217.930 131.985 ;
        RECT 218.120 131.815 218.290 131.985 ;
        RECT 218.480 131.815 218.650 131.985 ;
        RECT 218.840 131.815 219.010 131.985 ;
        RECT 219.200 131.815 219.370 131.985 ;
        RECT 219.560 131.815 219.730 131.985 ;
        RECT 219.920 131.815 220.090 131.985 ;
        RECT 220.280 131.815 220.450 131.985 ;
        RECT 220.640 131.815 220.810 131.985 ;
        RECT 221.000 131.815 221.170 131.985 ;
        RECT 221.360 131.815 221.530 131.985 ;
        RECT 221.720 131.815 221.890 131.985 ;
        RECT 222.080 131.815 222.250 131.985 ;
        RECT 222.440 131.815 222.610 131.985 ;
        RECT 222.800 131.815 222.970 131.985 ;
        RECT 223.160 131.815 223.330 131.985 ;
        RECT 223.520 131.815 223.690 131.985 ;
        RECT 223.880 131.815 224.050 131.985 ;
        RECT 224.240 131.815 224.410 131.985 ;
        RECT 224.600 131.815 224.770 131.985 ;
        RECT 224.960 131.815 225.130 131.985 ;
        RECT 225.320 131.815 225.490 131.985 ;
        RECT 225.680 131.815 225.850 131.985 ;
        RECT 226.040 131.815 226.210 131.985 ;
        RECT 226.400 131.815 226.570 131.985 ;
        RECT 226.760 131.815 226.930 131.985 ;
        RECT 227.120 131.815 227.290 131.985 ;
        RECT 227.480 131.815 227.650 131.985 ;
        RECT 227.840 131.815 228.010 131.985 ;
        RECT 228.200 131.815 228.370 131.985 ;
        RECT 228.560 131.815 228.730 131.985 ;
        RECT 228.920 131.815 229.090 131.985 ;
        RECT 258.020 131.300 258.190 131.470 ;
        RECT 258.380 131.300 258.550 131.470 ;
        RECT 258.740 131.300 258.910 131.470 ;
        RECT 259.100 131.300 259.270 131.470 ;
        RECT 259.460 131.300 259.630 131.470 ;
        RECT 259.820 131.300 259.990 131.470 ;
        RECT 260.180 131.300 260.350 131.470 ;
        RECT 260.540 131.300 260.710 131.470 ;
        RECT 260.900 131.300 261.070 131.470 ;
        RECT 261.260 131.300 261.430 131.470 ;
        RECT 261.620 131.300 261.790 131.470 ;
        RECT 261.980 131.300 262.150 131.470 ;
        RECT 262.340 131.300 262.510 131.470 ;
        RECT 262.700 131.300 262.870 131.470 ;
        RECT 263.060 131.300 263.230 131.470 ;
        RECT 263.420 131.300 263.590 131.470 ;
        RECT 263.780 131.300 263.950 131.470 ;
        RECT 264.140 131.300 264.310 131.470 ;
        RECT 264.500 131.300 264.670 131.470 ;
        RECT 264.860 131.300 265.030 131.470 ;
        RECT 265.220 131.300 265.390 131.470 ;
        RECT 265.580 131.300 265.750 131.470 ;
        RECT 265.940 131.300 266.110 131.470 ;
        RECT 266.300 131.300 266.470 131.470 ;
        RECT 266.660 131.300 266.830 131.470 ;
        RECT 267.020 131.300 267.190 131.470 ;
        RECT 267.380 131.300 267.550 131.470 ;
        RECT 267.740 131.300 267.910 131.470 ;
        RECT 268.100 131.300 268.270 131.470 ;
        RECT 268.460 131.300 268.630 131.470 ;
        RECT 268.820 131.300 268.990 131.470 ;
        RECT 269.180 131.300 269.350 131.470 ;
        RECT 269.540 131.300 269.710 131.470 ;
        RECT 269.900 131.300 270.070 131.470 ;
        RECT 270.260 131.300 270.430 131.470 ;
        RECT 270.620 131.300 270.790 131.470 ;
        RECT 270.980 131.300 271.150 131.470 ;
        RECT 271.340 131.300 271.510 131.470 ;
        RECT 271.700 131.300 271.870 131.470 ;
        RECT 272.060 131.300 272.230 131.470 ;
        RECT 272.420 131.300 272.590 131.470 ;
        RECT 272.780 131.300 272.950 131.470 ;
        RECT 273.140 131.300 273.310 131.470 ;
        RECT 273.500 131.300 273.670 131.470 ;
        RECT 273.860 131.300 274.030 131.470 ;
        RECT 274.220 131.300 274.390 131.470 ;
        RECT 274.580 131.300 274.750 131.470 ;
        RECT 274.940 131.300 275.110 131.470 ;
        RECT 275.300 131.300 275.470 131.470 ;
        RECT 275.660 131.300 275.830 131.470 ;
        RECT 276.020 131.300 276.190 131.470 ;
        RECT 276.380 131.300 276.550 131.470 ;
        RECT 276.740 131.300 276.910 131.470 ;
        RECT 277.100 131.300 277.270 131.470 ;
        RECT 277.460 131.300 277.630 131.470 ;
        RECT 277.820 131.300 277.990 131.470 ;
        RECT 278.180 131.300 278.350 131.470 ;
        RECT 271.770 98.050 272.300 98.580 ;
        RECT 275.455 99.340 275.625 99.510 ;
        RECT 275.455 98.980 275.625 99.150 ;
        RECT 275.455 98.620 275.625 98.790 ;
        RECT 273.290 98.390 273.460 98.560 ;
        RECT 275.455 98.260 275.625 98.430 ;
        RECT 275.455 97.900 275.625 98.070 ;
        RECT 275.455 97.540 275.625 97.710 ;
        RECT 275.455 97.180 275.625 97.350 ;
        RECT 275.455 96.820 275.625 96.990 ;
        RECT 275.455 96.460 275.625 96.630 ;
        RECT 275.455 96.100 275.625 96.270 ;
        RECT 271.765 95.195 272.295 95.725 ;
        RECT 273.290 95.610 273.460 95.780 ;
        RECT 275.455 95.740 275.625 95.910 ;
        RECT 275.455 95.380 275.625 95.550 ;
        RECT 275.455 95.020 275.625 95.190 ;
        RECT 275.455 94.660 275.625 94.830 ;
        RECT 271.765 92.445 272.295 92.975 ;
        RECT 273.290 92.830 273.460 93.000 ;
        RECT 275.090 92.685 275.620 93.215 ;
        RECT 276.920 92.820 277.090 92.990 ;
        RECT 275.070 90.715 275.600 91.245 ;
        RECT 276.920 90.830 277.090 91.000 ;
        RECT 271.750 89.665 272.280 90.195 ;
        RECT 273.290 90.050 273.460 90.220 ;
        RECT 258.660 88.760 258.830 88.930 ;
        RECT 258.660 88.400 258.830 88.570 ;
        RECT 258.660 88.040 258.830 88.210 ;
        RECT 258.660 87.680 258.830 87.850 ;
        RECT 209.575 83.845 209.745 84.015 ;
        RECT 209.935 83.845 210.105 84.015 ;
        RECT 210.295 83.845 210.465 84.015 ;
        RECT 210.655 83.845 210.825 84.015 ;
        RECT 211.015 83.845 211.185 84.015 ;
        RECT 211.375 83.845 211.545 84.015 ;
        RECT 211.735 83.845 211.905 84.015 ;
        RECT 212.095 83.845 212.265 84.015 ;
        RECT 212.455 83.845 212.625 84.015 ;
        RECT 212.815 83.845 212.985 84.015 ;
        RECT 213.175 83.845 213.345 84.015 ;
        RECT 213.535 83.845 213.705 84.015 ;
        RECT 213.895 83.845 214.065 84.015 ;
        RECT 214.255 83.845 214.425 84.015 ;
        RECT 214.615 83.845 214.785 84.015 ;
        RECT 214.975 83.845 215.145 84.015 ;
        RECT 215.335 83.845 215.505 84.015 ;
        RECT 215.695 83.845 215.865 84.015 ;
        RECT 216.055 83.845 216.225 84.015 ;
        RECT 216.415 83.845 216.585 84.015 ;
        RECT 216.775 83.845 216.945 84.015 ;
        RECT 217.135 83.845 217.305 84.015 ;
        RECT 217.495 83.845 217.665 84.015 ;
        RECT 217.855 83.845 218.025 84.015 ;
        RECT 218.215 83.845 218.385 84.015 ;
        RECT 218.575 83.845 218.745 84.015 ;
        RECT 218.935 83.845 219.105 84.015 ;
        RECT 219.295 83.845 219.465 84.015 ;
        RECT 219.655 83.845 219.825 84.015 ;
        RECT 220.015 83.845 220.185 84.015 ;
        RECT 220.375 83.845 220.545 84.015 ;
        RECT 220.735 83.845 220.905 84.015 ;
        RECT 221.095 83.845 221.265 84.015 ;
        RECT 221.455 83.845 221.625 84.015 ;
        RECT 221.815 83.845 221.985 84.015 ;
        RECT 222.175 83.845 222.345 84.015 ;
        RECT 222.535 83.845 222.705 84.015 ;
        RECT 222.895 83.845 223.065 84.015 ;
        RECT 223.255 83.845 223.425 84.015 ;
        RECT 223.615 83.845 223.785 84.015 ;
        RECT 223.975 83.845 224.145 84.015 ;
        RECT 224.335 83.845 224.505 84.015 ;
        RECT 224.695 83.845 224.865 84.015 ;
        RECT 225.055 83.845 225.225 84.015 ;
        RECT 225.415 83.845 225.585 84.015 ;
        RECT 225.775 83.845 225.945 84.015 ;
        RECT 226.135 83.845 226.305 84.015 ;
        RECT 226.495 83.845 226.665 84.015 ;
        RECT 226.855 83.845 227.025 84.015 ;
        RECT 227.215 83.845 227.385 84.015 ;
        RECT 227.575 83.845 227.745 84.015 ;
        RECT 227.935 83.845 228.105 84.015 ;
        RECT 228.295 83.845 228.465 84.015 ;
        RECT 228.655 83.845 228.825 84.015 ;
        RECT 229.015 83.845 229.185 84.015 ;
        RECT 259.260 86.200 259.430 86.370 ;
        RECT 259.260 85.840 259.430 86.010 ;
        RECT 259.260 85.480 259.430 85.650 ;
        RECT 259.260 85.120 259.430 85.290 ;
        RECT 259.260 84.760 259.430 84.930 ;
        RECT 259.260 84.400 259.430 84.570 ;
        RECT 259.260 84.040 259.430 84.210 ;
        RECT 259.260 83.680 259.430 83.850 ;
        RECT 271.750 86.875 272.280 87.405 ;
        RECT 273.290 87.270 273.460 87.440 ;
        RECT 275.130 86.950 275.660 87.480 ;
        RECT 276.920 87.260 277.090 87.430 ;
        RECT 271.765 84.380 272.295 84.910 ;
        RECT 273.290 84.490 273.460 84.660 ;
        RECT 209.575 82.330 209.745 82.500 ;
        RECT 209.935 82.330 210.105 82.500 ;
        RECT 210.295 82.330 210.465 82.500 ;
        RECT 210.655 82.330 210.825 82.500 ;
        RECT 211.015 82.330 211.185 82.500 ;
        RECT 211.375 82.330 211.545 82.500 ;
        RECT 211.735 82.330 211.905 82.500 ;
        RECT 212.095 82.330 212.265 82.500 ;
        RECT 212.455 82.330 212.625 82.500 ;
        RECT 212.815 82.330 212.985 82.500 ;
        RECT 213.175 82.330 213.345 82.500 ;
        RECT 213.535 82.330 213.705 82.500 ;
        RECT 213.895 82.330 214.065 82.500 ;
        RECT 214.255 82.330 214.425 82.500 ;
        RECT 214.615 82.330 214.785 82.500 ;
        RECT 214.975 82.330 215.145 82.500 ;
        RECT 215.335 82.330 215.505 82.500 ;
        RECT 215.695 82.330 215.865 82.500 ;
        RECT 216.055 82.330 216.225 82.500 ;
        RECT 216.415 82.330 216.585 82.500 ;
        RECT 216.775 82.330 216.945 82.500 ;
        RECT 217.135 82.330 217.305 82.500 ;
        RECT 217.495 82.330 217.665 82.500 ;
        RECT 217.855 82.330 218.025 82.500 ;
        RECT 218.215 82.330 218.385 82.500 ;
        RECT 218.575 82.330 218.745 82.500 ;
        RECT 218.935 82.330 219.105 82.500 ;
        RECT 219.295 82.330 219.465 82.500 ;
        RECT 219.655 82.330 219.825 82.500 ;
        RECT 220.015 82.330 220.185 82.500 ;
        RECT 220.375 82.330 220.545 82.500 ;
        RECT 220.735 82.330 220.905 82.500 ;
        RECT 221.095 82.330 221.265 82.500 ;
        RECT 221.455 82.330 221.625 82.500 ;
        RECT 221.815 82.330 221.985 82.500 ;
        RECT 222.175 82.330 222.345 82.500 ;
        RECT 222.535 82.330 222.705 82.500 ;
        RECT 222.895 82.330 223.065 82.500 ;
        RECT 223.255 82.330 223.425 82.500 ;
        RECT 223.615 82.330 223.785 82.500 ;
        RECT 223.975 82.330 224.145 82.500 ;
        RECT 224.335 82.330 224.505 82.500 ;
        RECT 224.695 82.330 224.865 82.500 ;
        RECT 225.055 82.330 225.225 82.500 ;
        RECT 225.415 82.330 225.585 82.500 ;
        RECT 225.775 82.330 225.945 82.500 ;
        RECT 226.135 82.330 226.305 82.500 ;
        RECT 226.495 82.330 226.665 82.500 ;
        RECT 226.855 82.330 227.025 82.500 ;
        RECT 227.215 82.330 227.385 82.500 ;
        RECT 227.575 82.330 227.745 82.500 ;
        RECT 227.935 82.330 228.105 82.500 ;
        RECT 228.295 82.330 228.465 82.500 ;
        RECT 228.655 82.330 228.825 82.500 ;
        RECT 229.015 82.330 229.185 82.500 ;
        RECT 258.225 79.295 258.395 79.465 ;
        RECT 258.225 78.935 258.395 79.105 ;
        RECT 259.835 79.090 260.005 79.260 ;
        RECT 258.225 78.575 258.395 78.745 ;
        RECT 258.225 78.215 258.395 78.385 ;
        RECT 258.310 76.825 259.200 77.715 ;
        RECT 258.215 76.115 258.385 76.285 ;
        RECT 258.215 75.755 258.385 75.925 ;
        RECT 258.215 75.395 258.385 75.565 ;
        RECT 259.825 75.270 259.995 75.440 ;
        RECT 258.215 75.035 258.385 75.205 ;
        RECT 279.645 79.295 279.815 79.465 ;
        RECT 278.035 79.090 278.205 79.260 ;
        RECT 279.645 78.935 279.815 79.105 ;
        RECT 279.645 78.575 279.815 78.745 ;
        RECT 279.645 78.215 279.815 78.385 ;
        RECT 278.840 76.825 279.730 77.715 ;
        RECT 279.655 76.115 279.825 76.285 ;
        RECT 279.655 75.755 279.825 75.925 ;
        RECT 278.045 75.270 278.215 75.440 ;
        RECT 279.655 75.395 279.825 75.565 ;
        RECT 279.655 75.035 279.825 75.205 ;
        RECT 209.550 65.905 209.720 66.075 ;
        RECT 209.910 65.905 210.080 66.075 ;
        RECT 210.270 65.905 210.440 66.075 ;
        RECT 210.630 65.905 210.800 66.075 ;
        RECT 210.990 65.905 211.160 66.075 ;
        RECT 211.350 65.905 211.520 66.075 ;
        RECT 211.710 65.905 211.880 66.075 ;
        RECT 212.070 65.905 212.240 66.075 ;
        RECT 212.430 65.905 212.600 66.075 ;
        RECT 212.790 65.905 212.960 66.075 ;
        RECT 213.150 65.905 213.320 66.075 ;
        RECT 213.510 65.905 213.680 66.075 ;
        RECT 213.870 65.905 214.040 66.075 ;
        RECT 214.230 65.905 214.400 66.075 ;
        RECT 214.590 65.905 214.760 66.075 ;
        RECT 214.950 65.905 215.120 66.075 ;
        RECT 215.310 65.905 215.480 66.075 ;
        RECT 215.670 65.905 215.840 66.075 ;
        RECT 216.030 65.905 216.200 66.075 ;
        RECT 216.390 65.905 216.560 66.075 ;
        RECT 216.750 65.905 216.920 66.075 ;
        RECT 217.110 65.905 217.280 66.075 ;
        RECT 217.470 65.905 217.640 66.075 ;
        RECT 217.830 65.905 218.000 66.075 ;
        RECT 218.190 65.905 218.360 66.075 ;
        RECT 218.550 65.905 218.720 66.075 ;
        RECT 218.910 65.905 219.080 66.075 ;
        RECT 219.270 65.905 219.440 66.075 ;
        RECT 219.630 65.905 219.800 66.075 ;
        RECT 219.990 65.905 220.160 66.075 ;
        RECT 220.350 65.905 220.520 66.075 ;
        RECT 220.710 65.905 220.880 66.075 ;
        RECT 221.070 65.905 221.240 66.075 ;
        RECT 221.430 65.905 221.600 66.075 ;
        RECT 221.790 65.905 221.960 66.075 ;
        RECT 222.150 65.905 222.320 66.075 ;
        RECT 222.510 65.905 222.680 66.075 ;
        RECT 222.870 65.905 223.040 66.075 ;
        RECT 223.230 65.905 223.400 66.075 ;
        RECT 223.590 65.905 223.760 66.075 ;
        RECT 223.950 65.905 224.120 66.075 ;
        RECT 224.310 65.905 224.480 66.075 ;
        RECT 224.670 65.905 224.840 66.075 ;
        RECT 225.030 65.905 225.200 66.075 ;
        RECT 225.390 65.905 225.560 66.075 ;
        RECT 225.750 65.905 225.920 66.075 ;
        RECT 226.110 65.905 226.280 66.075 ;
        RECT 226.470 65.905 226.640 66.075 ;
        RECT 226.830 65.905 227.000 66.075 ;
        RECT 227.190 65.905 227.360 66.075 ;
        RECT 227.550 65.905 227.720 66.075 ;
        RECT 227.910 65.905 228.080 66.075 ;
        RECT 228.270 65.905 228.440 66.075 ;
        RECT 228.630 65.905 228.800 66.075 ;
        RECT 228.990 65.905 229.160 66.075 ;
        RECT 286.730 65.815 286.900 65.985 ;
        RECT 287.090 65.815 287.260 65.985 ;
        RECT 287.450 65.815 287.620 65.985 ;
        RECT 287.810 65.815 287.980 65.985 ;
        RECT 288.170 65.815 288.340 65.985 ;
        RECT 288.530 65.815 288.700 65.985 ;
        RECT 288.890 65.815 289.060 65.985 ;
        RECT 289.250 65.815 289.420 65.985 ;
        RECT 289.610 65.815 289.780 65.985 ;
        RECT 289.970 65.815 290.140 65.985 ;
        RECT 290.330 65.815 290.500 65.985 ;
        RECT 290.690 65.815 290.860 65.985 ;
        RECT 291.050 65.815 291.220 65.985 ;
        RECT 291.410 65.815 291.580 65.985 ;
        RECT 291.770 65.815 291.940 65.985 ;
        RECT 292.130 65.815 292.300 65.985 ;
        RECT 292.490 65.815 292.660 65.985 ;
        RECT 292.850 65.815 293.020 65.985 ;
        RECT 293.210 65.815 293.380 65.985 ;
        RECT 293.570 65.815 293.740 65.985 ;
        RECT 293.930 65.815 294.100 65.985 ;
        RECT 294.290 65.815 294.460 65.985 ;
        RECT 294.650 65.815 294.820 65.985 ;
        RECT 295.010 65.815 295.180 65.985 ;
        RECT 295.370 65.815 295.540 65.985 ;
        RECT 295.730 65.815 295.900 65.985 ;
        RECT 296.090 65.815 296.260 65.985 ;
        RECT 296.450 65.815 296.620 65.985 ;
        RECT 296.810 65.815 296.980 65.985 ;
        RECT 297.170 65.815 297.340 65.985 ;
        RECT 297.530 65.815 297.700 65.985 ;
        RECT 297.890 65.815 298.060 65.985 ;
        RECT 298.250 65.815 298.420 65.985 ;
        RECT 298.610 65.815 298.780 65.985 ;
        RECT 298.970 65.815 299.140 65.985 ;
        RECT 299.330 65.815 299.500 65.985 ;
        RECT 299.690 65.815 299.860 65.985 ;
        RECT 300.050 65.815 300.220 65.985 ;
        RECT 300.410 65.815 300.580 65.985 ;
        RECT 300.770 65.815 300.940 65.985 ;
        RECT 301.130 65.815 301.300 65.985 ;
        RECT 301.490 65.815 301.660 65.985 ;
        RECT 301.850 65.815 302.020 65.985 ;
        RECT 302.210 65.815 302.380 65.985 ;
        RECT 302.570 65.815 302.740 65.985 ;
        RECT 302.930 65.815 303.100 65.985 ;
        RECT 303.290 65.815 303.460 65.985 ;
        RECT 303.650 65.815 303.820 65.985 ;
        RECT 304.010 65.815 304.180 65.985 ;
        RECT 304.370 65.815 304.540 65.985 ;
        RECT 304.730 65.815 304.900 65.985 ;
        RECT 305.090 65.815 305.260 65.985 ;
        RECT 305.450 65.815 305.620 65.985 ;
        RECT 305.810 65.815 305.980 65.985 ;
        RECT 306.170 65.815 306.340 65.985 ;
      LAYER met1 ;
        RECT 286.585 132.290 306.465 132.310 ;
        RECT 209.375 132.015 229.190 132.075 ;
        RECT 209.315 131.780 229.250 132.015 ;
        RECT 286.525 131.970 306.525 132.290 ;
        RECT 286.585 131.950 306.465 131.970 ;
        RECT 209.375 131.715 229.190 131.780 ;
        RECT 257.855 131.595 278.515 131.615 ;
        RECT 257.795 131.170 278.575 131.595 ;
        RECT 257.855 131.150 278.515 131.170 ;
        RECT 271.550 98.445 272.520 98.760 ;
        RECT 273.165 98.445 273.585 98.590 ;
        RECT 271.550 98.360 273.585 98.445 ;
        RECT 271.550 98.185 273.575 98.360 ;
        RECT 271.550 97.870 272.520 98.185 ;
        RECT 271.545 95.625 272.515 95.905 ;
        RECT 273.165 95.625 273.585 95.810 ;
        RECT 271.545 95.365 273.585 95.625 ;
        RECT 271.545 95.015 272.515 95.365 ;
        RECT 275.250 94.475 275.830 99.690 ;
        RECT 274.930 93.395 275.780 93.415 ;
        RECT 271.545 92.855 272.515 93.155 ;
        RECT 273.165 92.855 273.585 93.030 ;
        RECT 274.870 92.860 275.840 93.395 ;
        RECT 276.795 92.860 277.215 93.020 ;
        RECT 271.545 92.595 273.595 92.855 ;
        RECT 274.870 92.600 277.240 92.860 ;
        RECT 271.545 92.265 272.515 92.595 ;
        RECT 274.870 92.505 275.840 92.600 ;
        RECT 274.930 92.485 275.780 92.505 ;
        RECT 274.910 91.425 275.760 91.445 ;
        RECT 274.850 91.195 275.820 91.425 ;
        RECT 274.850 90.935 277.230 91.195 ;
        RECT 274.850 90.535 275.820 90.935 ;
        RECT 276.795 90.800 277.215 90.935 ;
        RECT 274.910 90.515 275.760 90.535 ;
        RECT 271.530 90.085 272.500 90.375 ;
        RECT 273.165 90.085 273.585 90.250 ;
        RECT 271.530 89.825 273.605 90.085 ;
        RECT 271.530 89.485 272.500 89.825 ;
        RECT 258.470 88.985 259.020 89.090 ;
        RECT 258.470 87.680 261.155 88.985 ;
        RECT 258.470 87.520 259.020 87.680 ;
        RECT 259.145 86.050 259.545 86.505 ;
        RECT 260.065 86.050 261.150 87.680 ;
        RECT 274.970 87.660 275.820 87.680 ;
        RECT 271.530 87.280 272.500 87.585 ;
        RECT 273.165 87.280 273.585 87.470 ;
        RECT 271.530 87.240 273.585 87.280 ;
        RECT 274.910 87.370 275.880 87.660 ;
        RECT 276.795 87.370 277.215 87.460 ;
        RECT 271.530 87.020 273.560 87.240 ;
        RECT 274.910 87.110 277.220 87.370 ;
        RECT 271.530 86.695 272.500 87.020 ;
        RECT 274.910 86.770 275.880 87.110 ;
        RECT 274.970 86.750 275.820 86.770 ;
        RECT 259.145 84.265 261.150 86.050 ;
        RECT 271.545 84.535 272.515 85.090 ;
        RECT 273.165 84.535 273.585 84.690 ;
        RECT 259.145 84.180 261.155 84.265 ;
        RECT 271.545 84.235 273.595 84.535 ;
        RECT 271.545 84.200 272.515 84.235 ;
        RECT 209.470 84.090 229.285 84.110 ;
        RECT 209.410 83.770 229.345 84.090 ;
        RECT 209.470 83.750 229.285 83.770 ;
        RECT 259.145 83.545 259.545 84.180 ;
        RECT 260.065 83.825 261.155 84.180 ;
        RECT 209.470 82.575 229.285 82.595 ;
        RECT 209.410 82.255 229.345 82.575 ;
        RECT 209.470 82.235 229.285 82.255 ;
        RECT 267.000 81.565 267.990 81.585 ;
        RECT 256.880 79.580 257.880 81.505 ;
        RECT 266.975 80.595 271.120 81.565 ;
        RECT 267.000 80.575 267.990 80.595 ;
        RECT 270.115 80.565 271.075 80.595 ;
        RECT 280.160 79.580 281.160 81.505 ;
        RECT 256.880 79.160 260.140 79.580 ;
        RECT 277.900 79.160 281.160 79.580 ;
        RECT 256.880 78.050 258.970 79.160 ;
        RECT 259.710 79.060 260.130 79.160 ;
        RECT 277.910 79.060 278.330 79.160 ;
        RECT 279.070 78.050 281.160 79.160 ;
        RECT 256.880 76.500 259.340 78.050 ;
        RECT 278.700 76.500 281.160 78.050 ;
        RECT 256.880 75.340 258.970 76.500 ;
        RECT 259.700 75.340 260.120 75.470 ;
        RECT 277.920 75.340 278.340 75.470 ;
        RECT 279.070 75.340 281.160 76.500 ;
        RECT 256.880 74.920 260.130 75.340 ;
        RECT 277.910 74.920 281.160 75.340 ;
        RECT 256.880 74.065 257.880 74.920 ;
        RECT 280.160 74.065 281.160 74.920 ;
        RECT 209.445 66.150 229.260 66.170 ;
        RECT 209.385 65.830 229.320 66.150 ;
        RECT 286.595 66.060 306.475 66.080 ;
        RECT 209.445 65.810 229.260 65.830 ;
        RECT 286.535 65.740 306.535 66.060 ;
        RECT 286.595 65.720 306.475 65.740 ;
      LAYER via ;
        RECT 209.395 131.765 209.655 132.025 ;
        RECT 209.715 131.765 209.975 132.025 ;
        RECT 210.035 131.765 210.295 132.025 ;
        RECT 210.355 131.765 210.615 132.025 ;
        RECT 210.675 131.765 210.935 132.025 ;
        RECT 210.995 131.765 211.255 132.025 ;
        RECT 211.315 131.765 211.575 132.025 ;
        RECT 211.635 131.765 211.895 132.025 ;
        RECT 211.955 131.765 212.215 132.025 ;
        RECT 212.275 131.765 212.535 132.025 ;
        RECT 212.595 131.765 212.855 132.025 ;
        RECT 212.915 131.765 213.175 132.025 ;
        RECT 213.235 131.765 213.495 132.025 ;
        RECT 213.555 131.765 213.815 132.025 ;
        RECT 213.875 131.765 214.135 132.025 ;
        RECT 214.195 131.765 214.455 132.025 ;
        RECT 214.515 131.765 214.775 132.025 ;
        RECT 214.835 131.765 215.095 132.025 ;
        RECT 215.155 131.765 215.415 132.025 ;
        RECT 215.475 131.765 215.735 132.025 ;
        RECT 215.795 131.765 216.055 132.025 ;
        RECT 216.115 131.765 216.375 132.025 ;
        RECT 216.435 131.765 216.695 132.025 ;
        RECT 216.755 131.765 217.015 132.025 ;
        RECT 217.075 131.765 217.335 132.025 ;
        RECT 217.395 131.765 217.655 132.025 ;
        RECT 217.715 131.765 217.975 132.025 ;
        RECT 218.035 131.765 218.295 132.025 ;
        RECT 218.355 131.765 218.615 132.025 ;
        RECT 218.675 131.765 218.935 132.025 ;
        RECT 218.995 131.765 219.255 132.025 ;
        RECT 219.315 131.765 219.575 132.025 ;
        RECT 219.635 131.765 219.895 132.025 ;
        RECT 219.955 131.765 220.215 132.025 ;
        RECT 220.275 131.765 220.535 132.025 ;
        RECT 220.595 131.765 220.855 132.025 ;
        RECT 220.915 131.765 221.175 132.025 ;
        RECT 221.235 131.765 221.495 132.025 ;
        RECT 221.555 131.765 221.815 132.025 ;
        RECT 221.875 131.765 222.135 132.025 ;
        RECT 222.195 131.765 222.455 132.025 ;
        RECT 222.515 131.765 222.775 132.025 ;
        RECT 222.835 131.765 223.095 132.025 ;
        RECT 223.155 131.765 223.415 132.025 ;
        RECT 223.475 131.765 223.735 132.025 ;
        RECT 223.795 131.765 224.055 132.025 ;
        RECT 224.115 131.765 224.375 132.025 ;
        RECT 224.435 131.765 224.695 132.025 ;
        RECT 224.755 131.765 225.015 132.025 ;
        RECT 225.075 131.765 225.335 132.025 ;
        RECT 225.395 131.765 225.655 132.025 ;
        RECT 225.715 131.765 225.975 132.025 ;
        RECT 226.035 131.765 226.295 132.025 ;
        RECT 226.355 131.765 226.615 132.025 ;
        RECT 226.675 131.765 226.935 132.025 ;
        RECT 226.995 131.765 227.255 132.025 ;
        RECT 227.315 131.765 227.575 132.025 ;
        RECT 227.635 131.765 227.895 132.025 ;
        RECT 227.955 131.765 228.215 132.025 ;
        RECT 228.275 131.765 228.535 132.025 ;
        RECT 228.595 131.765 228.855 132.025 ;
        RECT 228.915 131.765 229.175 132.025 ;
        RECT 286.635 132.000 286.895 132.260 ;
        RECT 286.955 132.000 287.215 132.260 ;
        RECT 287.275 132.000 287.535 132.260 ;
        RECT 287.595 132.000 287.855 132.260 ;
        RECT 287.915 132.000 288.175 132.260 ;
        RECT 288.235 132.000 288.495 132.260 ;
        RECT 288.555 132.000 288.815 132.260 ;
        RECT 288.875 132.000 289.135 132.260 ;
        RECT 289.195 132.000 289.455 132.260 ;
        RECT 289.515 132.000 289.775 132.260 ;
        RECT 289.835 132.000 290.095 132.260 ;
        RECT 290.155 132.000 290.415 132.260 ;
        RECT 290.475 132.000 290.735 132.260 ;
        RECT 290.795 132.000 291.055 132.260 ;
        RECT 291.115 132.000 291.375 132.260 ;
        RECT 291.435 132.000 291.695 132.260 ;
        RECT 291.755 132.000 292.015 132.260 ;
        RECT 292.075 132.000 292.335 132.260 ;
        RECT 292.395 132.000 292.655 132.260 ;
        RECT 292.715 132.000 292.975 132.260 ;
        RECT 293.035 132.000 293.295 132.260 ;
        RECT 293.355 132.000 293.615 132.260 ;
        RECT 293.675 132.000 293.935 132.260 ;
        RECT 293.995 132.000 294.255 132.260 ;
        RECT 294.315 132.000 294.575 132.260 ;
        RECT 294.635 132.000 294.895 132.260 ;
        RECT 294.955 132.000 295.215 132.260 ;
        RECT 295.275 132.000 295.535 132.260 ;
        RECT 295.595 132.000 295.855 132.260 ;
        RECT 295.915 132.000 296.175 132.260 ;
        RECT 296.235 132.000 296.495 132.260 ;
        RECT 296.555 132.000 296.815 132.260 ;
        RECT 296.875 132.000 297.135 132.260 ;
        RECT 297.195 132.000 297.455 132.260 ;
        RECT 297.515 132.000 297.775 132.260 ;
        RECT 297.835 132.000 298.095 132.260 ;
        RECT 298.155 132.000 298.415 132.260 ;
        RECT 298.475 132.000 298.735 132.260 ;
        RECT 298.795 132.000 299.055 132.260 ;
        RECT 299.115 132.000 299.375 132.260 ;
        RECT 299.435 132.000 299.695 132.260 ;
        RECT 299.755 132.000 300.015 132.260 ;
        RECT 300.075 132.000 300.335 132.260 ;
        RECT 300.395 132.000 300.655 132.260 ;
        RECT 300.715 132.000 300.975 132.260 ;
        RECT 301.035 132.000 301.295 132.260 ;
        RECT 301.355 132.000 301.615 132.260 ;
        RECT 301.675 132.000 301.935 132.260 ;
        RECT 301.995 132.000 302.255 132.260 ;
        RECT 302.315 132.000 302.575 132.260 ;
        RECT 302.635 132.000 302.895 132.260 ;
        RECT 302.955 132.000 303.215 132.260 ;
        RECT 303.275 132.000 303.535 132.260 ;
        RECT 303.595 132.000 303.855 132.260 ;
        RECT 303.915 132.000 304.175 132.260 ;
        RECT 304.235 132.000 304.495 132.260 ;
        RECT 304.555 132.000 304.815 132.260 ;
        RECT 304.875 132.000 305.135 132.260 ;
        RECT 305.195 132.000 305.455 132.260 ;
        RECT 305.515 132.000 305.775 132.260 ;
        RECT 305.835 132.000 306.095 132.260 ;
        RECT 306.155 132.000 306.415 132.260 ;
        RECT 257.975 131.255 258.235 131.515 ;
        RECT 258.295 131.255 258.555 131.515 ;
        RECT 258.615 131.255 258.875 131.515 ;
        RECT 258.935 131.255 259.195 131.515 ;
        RECT 259.255 131.255 259.515 131.515 ;
        RECT 259.575 131.255 259.835 131.515 ;
        RECT 259.895 131.255 260.155 131.515 ;
        RECT 260.215 131.255 260.475 131.515 ;
        RECT 260.535 131.255 260.795 131.515 ;
        RECT 260.855 131.255 261.115 131.515 ;
        RECT 261.175 131.255 261.435 131.515 ;
        RECT 261.495 131.255 261.755 131.515 ;
        RECT 261.815 131.255 262.075 131.515 ;
        RECT 262.135 131.255 262.395 131.515 ;
        RECT 262.455 131.255 262.715 131.515 ;
        RECT 262.775 131.255 263.035 131.515 ;
        RECT 263.095 131.255 263.355 131.515 ;
        RECT 263.415 131.255 263.675 131.515 ;
        RECT 263.735 131.255 263.995 131.515 ;
        RECT 264.055 131.255 264.315 131.515 ;
        RECT 264.375 131.255 264.635 131.515 ;
        RECT 264.695 131.255 264.955 131.515 ;
        RECT 265.015 131.255 265.275 131.515 ;
        RECT 265.335 131.255 265.595 131.515 ;
        RECT 265.655 131.255 265.915 131.515 ;
        RECT 265.975 131.255 266.235 131.515 ;
        RECT 266.295 131.255 266.555 131.515 ;
        RECT 266.615 131.255 266.875 131.515 ;
        RECT 266.935 131.255 267.195 131.515 ;
        RECT 267.255 131.255 267.515 131.515 ;
        RECT 267.575 131.255 267.835 131.515 ;
        RECT 267.895 131.255 268.155 131.515 ;
        RECT 268.215 131.255 268.475 131.515 ;
        RECT 268.535 131.255 268.795 131.515 ;
        RECT 268.855 131.255 269.115 131.515 ;
        RECT 269.175 131.255 269.435 131.515 ;
        RECT 269.495 131.255 269.755 131.515 ;
        RECT 269.815 131.255 270.075 131.515 ;
        RECT 270.135 131.255 270.395 131.515 ;
        RECT 270.455 131.255 270.715 131.515 ;
        RECT 270.775 131.255 271.035 131.515 ;
        RECT 271.095 131.255 271.355 131.515 ;
        RECT 271.415 131.255 271.675 131.515 ;
        RECT 271.735 131.255 271.995 131.515 ;
        RECT 272.055 131.255 272.315 131.515 ;
        RECT 272.375 131.255 272.635 131.515 ;
        RECT 272.695 131.255 272.955 131.515 ;
        RECT 273.015 131.255 273.275 131.515 ;
        RECT 273.335 131.255 273.595 131.515 ;
        RECT 273.655 131.255 273.915 131.515 ;
        RECT 273.975 131.255 274.235 131.515 ;
        RECT 274.295 131.255 274.555 131.515 ;
        RECT 274.615 131.255 274.875 131.515 ;
        RECT 274.935 131.255 275.195 131.515 ;
        RECT 275.255 131.255 275.515 131.515 ;
        RECT 275.575 131.255 275.835 131.515 ;
        RECT 275.895 131.255 276.155 131.515 ;
        RECT 276.215 131.255 276.475 131.515 ;
        RECT 276.535 131.255 276.795 131.515 ;
        RECT 276.855 131.255 277.115 131.515 ;
        RECT 277.175 131.255 277.435 131.515 ;
        RECT 277.495 131.255 277.755 131.515 ;
        RECT 277.815 131.255 278.075 131.515 ;
        RECT 278.135 131.255 278.395 131.515 ;
        RECT 275.410 99.355 275.670 99.615 ;
        RECT 275.410 99.035 275.670 99.295 ;
        RECT 275.410 98.715 275.670 98.975 ;
        RECT 275.410 98.395 275.670 98.655 ;
        RECT 275.410 98.075 275.670 98.335 ;
        RECT 275.410 97.755 275.670 98.015 ;
        RECT 275.410 97.435 275.670 97.695 ;
        RECT 275.410 97.115 275.670 97.375 ;
        RECT 275.410 96.795 275.670 97.055 ;
        RECT 275.410 96.475 275.670 96.735 ;
        RECT 275.410 96.155 275.670 96.415 ;
        RECT 275.410 95.835 275.670 96.095 ;
        RECT 275.410 95.515 275.670 95.775 ;
        RECT 275.410 95.195 275.670 95.455 ;
        RECT 275.410 94.875 275.670 95.135 ;
        RECT 275.410 94.555 275.670 94.815 ;
        RECT 275.065 92.660 275.645 93.240 ;
        RECT 275.045 90.690 275.625 91.270 ;
        RECT 275.105 86.925 275.685 87.505 ;
        RECT 209.490 83.800 209.750 84.060 ;
        RECT 209.810 83.800 210.070 84.060 ;
        RECT 210.130 83.800 210.390 84.060 ;
        RECT 210.450 83.800 210.710 84.060 ;
        RECT 210.770 83.800 211.030 84.060 ;
        RECT 211.090 83.800 211.350 84.060 ;
        RECT 211.410 83.800 211.670 84.060 ;
        RECT 211.730 83.800 211.990 84.060 ;
        RECT 212.050 83.800 212.310 84.060 ;
        RECT 212.370 83.800 212.630 84.060 ;
        RECT 212.690 83.800 212.950 84.060 ;
        RECT 213.010 83.800 213.270 84.060 ;
        RECT 213.330 83.800 213.590 84.060 ;
        RECT 213.650 83.800 213.910 84.060 ;
        RECT 213.970 83.800 214.230 84.060 ;
        RECT 214.290 83.800 214.550 84.060 ;
        RECT 214.610 83.800 214.870 84.060 ;
        RECT 214.930 83.800 215.190 84.060 ;
        RECT 215.250 83.800 215.510 84.060 ;
        RECT 215.570 83.800 215.830 84.060 ;
        RECT 215.890 83.800 216.150 84.060 ;
        RECT 216.210 83.800 216.470 84.060 ;
        RECT 216.530 83.800 216.790 84.060 ;
        RECT 216.850 83.800 217.110 84.060 ;
        RECT 217.170 83.800 217.430 84.060 ;
        RECT 217.490 83.800 217.750 84.060 ;
        RECT 217.810 83.800 218.070 84.060 ;
        RECT 218.130 83.800 218.390 84.060 ;
        RECT 218.450 83.800 218.710 84.060 ;
        RECT 218.770 83.800 219.030 84.060 ;
        RECT 219.090 83.800 219.350 84.060 ;
        RECT 219.410 83.800 219.670 84.060 ;
        RECT 219.730 83.800 219.990 84.060 ;
        RECT 220.050 83.800 220.310 84.060 ;
        RECT 220.370 83.800 220.630 84.060 ;
        RECT 220.690 83.800 220.950 84.060 ;
        RECT 221.010 83.800 221.270 84.060 ;
        RECT 221.330 83.800 221.590 84.060 ;
        RECT 221.650 83.800 221.910 84.060 ;
        RECT 221.970 83.800 222.230 84.060 ;
        RECT 222.290 83.800 222.550 84.060 ;
        RECT 222.610 83.800 222.870 84.060 ;
        RECT 222.930 83.800 223.190 84.060 ;
        RECT 223.250 83.800 223.510 84.060 ;
        RECT 223.570 83.800 223.830 84.060 ;
        RECT 223.890 83.800 224.150 84.060 ;
        RECT 224.210 83.800 224.470 84.060 ;
        RECT 224.530 83.800 224.790 84.060 ;
        RECT 224.850 83.800 225.110 84.060 ;
        RECT 225.170 83.800 225.430 84.060 ;
        RECT 225.490 83.800 225.750 84.060 ;
        RECT 225.810 83.800 226.070 84.060 ;
        RECT 226.130 83.800 226.390 84.060 ;
        RECT 226.450 83.800 226.710 84.060 ;
        RECT 226.770 83.800 227.030 84.060 ;
        RECT 227.090 83.800 227.350 84.060 ;
        RECT 227.410 83.800 227.670 84.060 ;
        RECT 227.730 83.800 227.990 84.060 ;
        RECT 228.050 83.800 228.310 84.060 ;
        RECT 228.370 83.800 228.630 84.060 ;
        RECT 228.690 83.800 228.950 84.060 ;
        RECT 229.010 83.800 229.270 84.060 ;
        RECT 260.160 83.915 260.420 84.175 ;
        RECT 260.480 83.915 260.740 84.175 ;
        RECT 260.800 83.915 261.060 84.175 ;
        RECT 209.490 82.285 209.750 82.545 ;
        RECT 209.810 82.285 210.070 82.545 ;
        RECT 210.130 82.285 210.390 82.545 ;
        RECT 210.450 82.285 210.710 82.545 ;
        RECT 210.770 82.285 211.030 82.545 ;
        RECT 211.090 82.285 211.350 82.545 ;
        RECT 211.410 82.285 211.670 82.545 ;
        RECT 211.730 82.285 211.990 82.545 ;
        RECT 212.050 82.285 212.310 82.545 ;
        RECT 212.370 82.285 212.630 82.545 ;
        RECT 212.690 82.285 212.950 82.545 ;
        RECT 213.010 82.285 213.270 82.545 ;
        RECT 213.330 82.285 213.590 82.545 ;
        RECT 213.650 82.285 213.910 82.545 ;
        RECT 213.970 82.285 214.230 82.545 ;
        RECT 214.290 82.285 214.550 82.545 ;
        RECT 214.610 82.285 214.870 82.545 ;
        RECT 214.930 82.285 215.190 82.545 ;
        RECT 215.250 82.285 215.510 82.545 ;
        RECT 215.570 82.285 215.830 82.545 ;
        RECT 215.890 82.285 216.150 82.545 ;
        RECT 216.210 82.285 216.470 82.545 ;
        RECT 216.530 82.285 216.790 82.545 ;
        RECT 216.850 82.285 217.110 82.545 ;
        RECT 217.170 82.285 217.430 82.545 ;
        RECT 217.490 82.285 217.750 82.545 ;
        RECT 217.810 82.285 218.070 82.545 ;
        RECT 218.130 82.285 218.390 82.545 ;
        RECT 218.450 82.285 218.710 82.545 ;
        RECT 218.770 82.285 219.030 82.545 ;
        RECT 219.090 82.285 219.350 82.545 ;
        RECT 219.410 82.285 219.670 82.545 ;
        RECT 219.730 82.285 219.990 82.545 ;
        RECT 220.050 82.285 220.310 82.545 ;
        RECT 220.370 82.285 220.630 82.545 ;
        RECT 220.690 82.285 220.950 82.545 ;
        RECT 221.010 82.285 221.270 82.545 ;
        RECT 221.330 82.285 221.590 82.545 ;
        RECT 221.650 82.285 221.910 82.545 ;
        RECT 221.970 82.285 222.230 82.545 ;
        RECT 222.290 82.285 222.550 82.545 ;
        RECT 222.610 82.285 222.870 82.545 ;
        RECT 222.930 82.285 223.190 82.545 ;
        RECT 223.250 82.285 223.510 82.545 ;
        RECT 223.570 82.285 223.830 82.545 ;
        RECT 223.890 82.285 224.150 82.545 ;
        RECT 224.210 82.285 224.470 82.545 ;
        RECT 224.530 82.285 224.790 82.545 ;
        RECT 224.850 82.285 225.110 82.545 ;
        RECT 225.170 82.285 225.430 82.545 ;
        RECT 225.490 82.285 225.750 82.545 ;
        RECT 225.810 82.285 226.070 82.545 ;
        RECT 226.130 82.285 226.390 82.545 ;
        RECT 226.450 82.285 226.710 82.545 ;
        RECT 226.770 82.285 227.030 82.545 ;
        RECT 227.090 82.285 227.350 82.545 ;
        RECT 227.410 82.285 227.670 82.545 ;
        RECT 227.730 82.285 227.990 82.545 ;
        RECT 228.050 82.285 228.310 82.545 ;
        RECT 228.370 82.285 228.630 82.545 ;
        RECT 228.690 82.285 228.950 82.545 ;
        RECT 229.010 82.285 229.270 82.545 ;
        RECT 257.150 74.265 257.730 81.245 ;
        RECT 267.045 80.630 267.945 81.530 ;
        RECT 270.145 80.775 271.045 81.355 ;
        RECT 280.440 74.275 281.020 81.255 ;
        RECT 209.465 65.860 209.725 66.120 ;
        RECT 209.785 65.860 210.045 66.120 ;
        RECT 210.105 65.860 210.365 66.120 ;
        RECT 210.425 65.860 210.685 66.120 ;
        RECT 210.745 65.860 211.005 66.120 ;
        RECT 211.065 65.860 211.325 66.120 ;
        RECT 211.385 65.860 211.645 66.120 ;
        RECT 211.705 65.860 211.965 66.120 ;
        RECT 212.025 65.860 212.285 66.120 ;
        RECT 212.345 65.860 212.605 66.120 ;
        RECT 212.665 65.860 212.925 66.120 ;
        RECT 212.985 65.860 213.245 66.120 ;
        RECT 213.305 65.860 213.565 66.120 ;
        RECT 213.625 65.860 213.885 66.120 ;
        RECT 213.945 65.860 214.205 66.120 ;
        RECT 214.265 65.860 214.525 66.120 ;
        RECT 214.585 65.860 214.845 66.120 ;
        RECT 214.905 65.860 215.165 66.120 ;
        RECT 215.225 65.860 215.485 66.120 ;
        RECT 215.545 65.860 215.805 66.120 ;
        RECT 215.865 65.860 216.125 66.120 ;
        RECT 216.185 65.860 216.445 66.120 ;
        RECT 216.505 65.860 216.765 66.120 ;
        RECT 216.825 65.860 217.085 66.120 ;
        RECT 217.145 65.860 217.405 66.120 ;
        RECT 217.465 65.860 217.725 66.120 ;
        RECT 217.785 65.860 218.045 66.120 ;
        RECT 218.105 65.860 218.365 66.120 ;
        RECT 218.425 65.860 218.685 66.120 ;
        RECT 218.745 65.860 219.005 66.120 ;
        RECT 219.065 65.860 219.325 66.120 ;
        RECT 219.385 65.860 219.645 66.120 ;
        RECT 219.705 65.860 219.965 66.120 ;
        RECT 220.025 65.860 220.285 66.120 ;
        RECT 220.345 65.860 220.605 66.120 ;
        RECT 220.665 65.860 220.925 66.120 ;
        RECT 220.985 65.860 221.245 66.120 ;
        RECT 221.305 65.860 221.565 66.120 ;
        RECT 221.625 65.860 221.885 66.120 ;
        RECT 221.945 65.860 222.205 66.120 ;
        RECT 222.265 65.860 222.525 66.120 ;
        RECT 222.585 65.860 222.845 66.120 ;
        RECT 222.905 65.860 223.165 66.120 ;
        RECT 223.225 65.860 223.485 66.120 ;
        RECT 223.545 65.860 223.805 66.120 ;
        RECT 223.865 65.860 224.125 66.120 ;
        RECT 224.185 65.860 224.445 66.120 ;
        RECT 224.505 65.860 224.765 66.120 ;
        RECT 224.825 65.860 225.085 66.120 ;
        RECT 225.145 65.860 225.405 66.120 ;
        RECT 225.465 65.860 225.725 66.120 ;
        RECT 225.785 65.860 226.045 66.120 ;
        RECT 226.105 65.860 226.365 66.120 ;
        RECT 226.425 65.860 226.685 66.120 ;
        RECT 226.745 65.860 227.005 66.120 ;
        RECT 227.065 65.860 227.325 66.120 ;
        RECT 227.385 65.860 227.645 66.120 ;
        RECT 227.705 65.860 227.965 66.120 ;
        RECT 228.025 65.860 228.285 66.120 ;
        RECT 228.345 65.860 228.605 66.120 ;
        RECT 228.665 65.860 228.925 66.120 ;
        RECT 228.985 65.860 229.245 66.120 ;
        RECT 286.645 65.770 286.905 66.030 ;
        RECT 286.965 65.770 287.225 66.030 ;
        RECT 287.285 65.770 287.545 66.030 ;
        RECT 287.605 65.770 287.865 66.030 ;
        RECT 287.925 65.770 288.185 66.030 ;
        RECT 288.245 65.770 288.505 66.030 ;
        RECT 288.565 65.770 288.825 66.030 ;
        RECT 288.885 65.770 289.145 66.030 ;
        RECT 289.205 65.770 289.465 66.030 ;
        RECT 289.525 65.770 289.785 66.030 ;
        RECT 289.845 65.770 290.105 66.030 ;
        RECT 290.165 65.770 290.425 66.030 ;
        RECT 290.485 65.770 290.745 66.030 ;
        RECT 290.805 65.770 291.065 66.030 ;
        RECT 291.125 65.770 291.385 66.030 ;
        RECT 291.445 65.770 291.705 66.030 ;
        RECT 291.765 65.770 292.025 66.030 ;
        RECT 292.085 65.770 292.345 66.030 ;
        RECT 292.405 65.770 292.665 66.030 ;
        RECT 292.725 65.770 292.985 66.030 ;
        RECT 293.045 65.770 293.305 66.030 ;
        RECT 293.365 65.770 293.625 66.030 ;
        RECT 293.685 65.770 293.945 66.030 ;
        RECT 294.005 65.770 294.265 66.030 ;
        RECT 294.325 65.770 294.585 66.030 ;
        RECT 294.645 65.770 294.905 66.030 ;
        RECT 294.965 65.770 295.225 66.030 ;
        RECT 295.285 65.770 295.545 66.030 ;
        RECT 295.605 65.770 295.865 66.030 ;
        RECT 295.925 65.770 296.185 66.030 ;
        RECT 296.245 65.770 296.505 66.030 ;
        RECT 296.565 65.770 296.825 66.030 ;
        RECT 296.885 65.770 297.145 66.030 ;
        RECT 297.205 65.770 297.465 66.030 ;
        RECT 297.525 65.770 297.785 66.030 ;
        RECT 297.845 65.770 298.105 66.030 ;
        RECT 298.165 65.770 298.425 66.030 ;
        RECT 298.485 65.770 298.745 66.030 ;
        RECT 298.805 65.770 299.065 66.030 ;
        RECT 299.125 65.770 299.385 66.030 ;
        RECT 299.445 65.770 299.705 66.030 ;
        RECT 299.765 65.770 300.025 66.030 ;
        RECT 300.085 65.770 300.345 66.030 ;
        RECT 300.405 65.770 300.665 66.030 ;
        RECT 300.725 65.770 300.985 66.030 ;
        RECT 301.045 65.770 301.305 66.030 ;
        RECT 301.365 65.770 301.625 66.030 ;
        RECT 301.685 65.770 301.945 66.030 ;
        RECT 302.005 65.770 302.265 66.030 ;
        RECT 302.325 65.770 302.585 66.030 ;
        RECT 302.645 65.770 302.905 66.030 ;
        RECT 302.965 65.770 303.225 66.030 ;
        RECT 303.285 65.770 303.545 66.030 ;
        RECT 303.605 65.770 303.865 66.030 ;
        RECT 303.925 65.770 304.185 66.030 ;
        RECT 304.245 65.770 304.505 66.030 ;
        RECT 304.565 65.770 304.825 66.030 ;
        RECT 304.885 65.770 305.145 66.030 ;
        RECT 305.205 65.770 305.465 66.030 ;
        RECT 305.525 65.770 305.785 66.030 ;
        RECT 305.845 65.770 306.105 66.030 ;
        RECT 306.165 65.770 306.425 66.030 ;
      LAYER met2 ;
        RECT 209.330 132.025 229.330 134.100 ;
        RECT 209.325 131.765 229.330 132.025 ;
        RECT 286.515 131.985 306.515 134.100 ;
        RECT 209.330 84.060 229.330 131.765 ;
        RECT 257.215 130.965 306.515 131.985 ;
        RECT 260.160 103.085 277.720 130.965 ;
        RECT 286.515 100.815 306.515 130.965 ;
        RECT 274.745 94.785 306.515 100.815 ;
        RECT 274.745 90.260 279.875 94.785 ;
        RECT 277.110 89.950 279.875 90.260 ;
        RECT 286.515 89.950 306.515 94.785 ;
        RECT 277.110 88.535 306.515 89.950 ;
        RECT 274.760 86.555 306.515 88.535 ;
        RECT 209.330 83.800 229.335 84.060 ;
        RECT 260.015 83.875 261.205 84.215 ;
        RECT 280.540 83.920 306.515 86.555 ;
        RECT 209.330 82.545 229.330 83.800 ;
        RECT 209.330 82.285 229.335 82.545 ;
        RECT 209.330 63.930 229.330 82.285 ;
        RECT 260.065 81.530 261.150 83.875 ;
        RECT 266.950 81.530 268.040 81.535 ;
        RECT 254.865 80.625 268.040 81.530 ;
        RECT 270.065 81.475 271.125 81.510 ;
        RECT 286.515 81.475 306.515 83.920 ;
        RECT 254.865 80.550 267.995 80.625 ;
        RECT 270.065 80.615 306.515 81.475 ;
        RECT 270.110 80.590 306.515 80.615 ;
        RECT 254.865 74.075 257.895 80.550 ;
        RECT 280.140 74.050 306.515 80.590 ;
        RECT 286.515 66.030 306.515 74.050 ;
        RECT 286.515 65.770 306.525 66.030 ;
        RECT 286.515 63.930 306.515 65.770 ;
      LAYER via2 ;
        RECT 214.575 132.565 216.055 134.000 ;
        RECT 217.905 132.565 219.385 134.000 ;
        RECT 221.200 132.545 222.680 133.980 ;
        RECT 224.515 132.545 225.995 133.980 ;
        RECT 291.760 132.565 293.240 134.000 ;
        RECT 295.090 132.565 296.570 134.000 ;
        RECT 298.385 132.545 299.865 133.980 ;
        RECT 301.700 132.545 303.180 133.980 ;
        RECT 214.575 64.105 216.055 65.540 ;
        RECT 217.905 64.105 219.385 65.540 ;
        RECT 221.200 64.085 222.680 65.520 ;
        RECT 224.515 64.085 225.995 65.520 ;
        RECT 291.760 64.105 293.240 65.540 ;
        RECT 295.090 64.105 296.570 65.540 ;
        RECT 298.385 64.085 299.865 65.520 ;
        RECT 301.700 64.085 303.180 65.520 ;
      LAYER met3 ;
        RECT 209.330 132.390 229.330 134.100 ;
        RECT 286.515 132.390 306.515 134.100 ;
        RECT 209.330 63.930 229.330 65.640 ;
        RECT 286.515 63.930 306.515 65.640 ;
      LAYER via3 ;
        RECT 214.555 132.545 216.075 134.020 ;
        RECT 217.885 132.545 219.405 134.020 ;
        RECT 221.180 132.525 222.700 134.000 ;
        RECT 224.495 132.525 226.015 134.000 ;
        RECT 291.740 132.545 293.260 134.020 ;
        RECT 295.070 132.545 296.590 134.020 ;
        RECT 298.365 132.525 299.885 134.000 ;
        RECT 301.680 132.525 303.200 134.000 ;
        RECT 214.555 64.085 216.075 65.560 ;
        RECT 217.885 64.085 219.405 65.560 ;
        RECT 221.180 64.065 222.700 65.540 ;
        RECT 224.495 64.065 226.015 65.540 ;
        RECT 291.740 64.085 293.260 65.560 ;
        RECT 295.070 64.085 296.590 65.560 ;
        RECT 298.365 64.065 299.885 65.540 ;
        RECT 301.680 64.065 303.200 65.540 ;
      LAYER met4 ;
        RECT 214.545 3.300 216.145 211.800 ;
        RECT 217.845 3.300 219.445 211.800 ;
        RECT 221.145 3.300 222.745 211.800 ;
        RECT 224.445 3.300 226.045 211.800 ;
        RECT 291.730 3.300 293.330 211.800 ;
        RECT 295.030 3.300 296.630 211.800 ;
        RECT 298.330 3.300 299.930 211.800 ;
        RECT 301.630 3.300 303.230 211.800 ;
    END
  END vssa1
  PIN vssd1
    ANTENNADIFFAREA 15.428800 ;
    PORT
      LAYER pwell ;
        RECT 261.245 71.360 276.965 71.790 ;
        RECT 261.245 69.970 261.675 71.360 ;
        RECT 276.535 69.970 276.965 71.360 ;
        RECT 277.885 70.460 279.615 72.190 ;
        RECT 261.245 69.540 276.965 69.970 ;
        RECT 258.710 67.250 259.440 68.580 ;
        RECT 260.340 66.470 263.030 68.480 ;
        RECT 267.245 66.045 269.435 68.055 ;
        RECT 275.010 66.470 277.700 68.480 ;
        RECT 278.600 67.250 279.330 68.580 ;
        RECT 260.510 64.310 262.240 66.040 ;
        RECT 267.245 63.980 269.435 65.990 ;
        RECT 269.535 63.980 271.645 65.990 ;
      LAYER li1 ;
        RECT 278.015 71.890 279.485 72.060 ;
        RECT 261.375 71.490 276.835 71.660 ;
        RECT 261.375 69.840 261.545 71.490 ;
        RECT 276.665 69.840 276.835 71.490 ;
        RECT 261.375 69.670 276.835 69.840 ;
        RECT 278.015 70.760 278.185 71.890 ;
        RECT 279.315 70.760 279.485 71.890 ;
        RECT 278.015 70.590 279.485 70.760 ;
        RECT 261.375 69.140 276.825 69.670 ;
        RECT 278.015 68.980 279.030 70.590 ;
        RECT 260.150 68.410 262.900 68.560 ;
        RECT 258.840 68.180 262.900 68.410 ;
        RECT 258.840 67.060 260.660 68.180 ;
        RECT 261.010 67.170 262.050 67.340 ;
        RECT 260.150 66.770 260.660 67.060 ;
        RECT 262.730 66.770 262.900 68.180 ;
        RECT 275.140 68.410 277.890 68.560 ;
        RECT 275.140 68.180 279.200 68.410 ;
        RECT 269.310 67.925 269.660 67.930 ;
        RECT 260.150 66.600 262.900 66.770 ;
        RECT 267.375 67.755 269.675 67.925 ;
        RECT 260.150 66.570 262.105 66.600 ;
        RECT 260.190 65.910 262.105 66.570 ;
        RECT 267.375 66.345 267.545 67.755 ;
        RECT 268.225 67.185 268.765 67.355 ;
        RECT 269.135 66.345 269.675 67.755 ;
        RECT 275.140 66.770 275.310 68.180 ;
        RECT 275.990 67.170 277.030 67.340 ;
        RECT 277.380 67.060 279.200 68.180 ;
        RECT 277.380 66.770 277.890 67.060 ;
        RECT 275.140 66.600 277.890 66.770 ;
        RECT 277.380 66.570 277.890 66.600 ;
        RECT 267.375 66.175 269.675 66.345 ;
        RECT 260.190 65.740 262.110 65.910 ;
        RECT 267.380 65.860 269.675 66.175 ;
        RECT 260.190 64.610 260.810 65.740 ;
        RECT 261.940 64.610 262.110 65.740 ;
        RECT 260.190 64.445 262.110 64.610 ;
        RECT 260.640 64.440 262.110 64.445 ;
        RECT 267.375 65.690 271.515 65.860 ;
        RECT 267.375 64.280 267.545 65.690 ;
        RECT 269.135 64.280 269.835 65.690 ;
        RECT 270.515 65.120 270.975 65.290 ;
        RECT 271.345 64.280 271.515 65.690 ;
        RECT 267.375 64.110 271.515 64.280 ;
        RECT 269.300 64.060 269.675 64.110 ;
      LAYER mcon ;
        RECT 261.935 69.335 262.105 69.505 ;
        RECT 262.295 69.335 262.465 69.505 ;
        RECT 262.655 69.335 262.825 69.505 ;
        RECT 263.015 69.335 263.185 69.505 ;
        RECT 263.375 69.335 263.545 69.505 ;
        RECT 263.735 69.335 263.905 69.505 ;
        RECT 264.095 69.335 264.265 69.505 ;
        RECT 264.455 69.335 264.625 69.505 ;
        RECT 264.815 69.335 264.985 69.505 ;
        RECT 265.175 69.335 265.345 69.505 ;
        RECT 265.535 69.335 265.705 69.505 ;
        RECT 265.895 69.335 266.065 69.505 ;
        RECT 266.255 69.335 266.425 69.505 ;
        RECT 266.615 69.335 266.785 69.505 ;
        RECT 266.975 69.335 267.145 69.505 ;
        RECT 267.335 69.335 267.505 69.505 ;
        RECT 267.695 69.335 267.865 69.505 ;
        RECT 268.055 69.335 268.225 69.505 ;
        RECT 268.415 69.335 268.585 69.505 ;
        RECT 268.775 69.335 268.945 69.505 ;
        RECT 269.135 69.335 269.305 69.505 ;
        RECT 269.495 69.335 269.665 69.505 ;
        RECT 269.855 69.335 270.025 69.505 ;
        RECT 270.215 69.335 270.385 69.505 ;
        RECT 270.575 69.335 270.745 69.505 ;
        RECT 270.935 69.335 271.105 69.505 ;
        RECT 271.295 69.335 271.465 69.505 ;
        RECT 271.655 69.335 271.825 69.505 ;
        RECT 272.015 69.335 272.185 69.505 ;
        RECT 272.375 69.335 272.545 69.505 ;
        RECT 272.735 69.335 272.905 69.505 ;
        RECT 273.095 69.335 273.265 69.505 ;
        RECT 273.455 69.335 273.625 69.505 ;
        RECT 273.815 69.335 273.985 69.505 ;
        RECT 274.175 69.335 274.345 69.505 ;
        RECT 274.535 69.335 274.705 69.505 ;
        RECT 274.895 69.335 275.065 69.505 ;
        RECT 275.255 69.335 275.425 69.505 ;
        RECT 275.615 69.335 275.785 69.505 ;
        RECT 275.975 69.335 276.145 69.505 ;
        RECT 278.080 69.180 278.970 69.710 ;
        RECT 259.650 67.370 260.180 67.900 ;
        RECT 261.265 67.170 261.435 67.340 ;
        RECT 261.625 67.170 261.795 67.340 ;
        RECT 269.405 67.635 269.575 67.805 ;
        RECT 268.410 67.185 268.580 67.355 ;
        RECT 269.405 67.275 269.575 67.445 ;
        RECT 269.405 66.915 269.575 67.085 ;
        RECT 269.405 66.555 269.575 66.725 ;
        RECT 277.860 67.370 278.390 67.900 ;
        RECT 276.245 67.170 276.415 67.340 ;
        RECT 276.605 67.170 276.775 67.340 ;
        RECT 269.405 66.195 269.575 66.365 ;
        RECT 269.405 65.835 269.575 66.005 ;
        RECT 269.405 65.475 269.575 65.645 ;
        RECT 269.405 65.115 269.575 65.285 ;
        RECT 270.660 65.120 270.830 65.290 ;
      LAYER met1 ;
        RECT 259.615 68.810 279.030 69.910 ;
        RECT 259.615 68.500 260.625 68.810 ;
        RECT 259.570 67.160 260.625 68.500 ;
        RECT 268.260 68.370 270.975 68.810 ;
        RECT 277.870 68.500 279.030 68.810 ;
        RECT 268.260 67.385 268.720 68.370 ;
        RECT 259.570 67.150 260.630 67.160 ;
        RECT 261.030 67.150 262.030 67.370 ;
        RECT 268.245 67.155 268.745 67.385 ;
        RECT 259.570 66.920 262.040 67.150 ;
        RECT 259.570 66.260 260.625 66.920 ;
        RECT 269.305 65.010 269.685 68.370 ;
        RECT 270.540 65.320 270.975 68.370 ;
        RECT 276.010 67.150 277.010 67.370 ;
        RECT 277.470 67.160 279.030 68.500 ;
        RECT 277.410 67.150 279.030 67.160 ;
        RECT 276.000 66.920 279.030 67.150 ;
        RECT 277.470 66.270 279.030 66.920 ;
        RECT 277.470 66.260 278.470 66.270 ;
        RECT 270.535 65.100 270.975 65.320 ;
        RECT 270.535 65.090 270.955 65.100 ;
      LAYER via ;
        RECT 259.840 66.490 260.420 67.070 ;
      LAYER met2 ;
        RECT 259.625 63.930 260.625 68.590 ;
      LAYER via2 ;
        RECT 259.825 64.300 260.505 68.100 ;
      LAYER met3 ;
        RECT 259.625 63.930 260.625 68.590 ;
      LAYER via3 ;
        RECT 259.805 64.280 260.525 68.120 ;
      LAYER met4 ;
        RECT 259.335 3.300 260.935 211.800 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER nwell ;
        RECT 263.120 66.420 265.960 68.530 ;
        RECT 272.080 66.420 274.920 68.530 ;
        RECT 263.165 63.930 266.005 66.420 ;
      LAYER li1 ;
        RECT 266.165 97.910 266.625 98.080 ;
        RECT 263.300 68.180 266.140 68.570 ;
        RECT 263.300 66.770 263.470 68.180 ;
        RECT 265.610 67.840 266.140 68.180 ;
        RECT 271.900 68.180 274.740 68.570 ;
        RECT 271.900 67.840 272.430 68.180 ;
        RECT 264.200 67.170 265.240 67.340 ;
        RECT 265.610 67.050 266.600 67.840 ;
        RECT 271.440 67.050 272.430 67.840 ;
        RECT 272.800 67.170 273.840 67.340 ;
        RECT 265.610 66.770 266.140 67.050 ;
        RECT 263.300 66.600 266.140 66.770 ;
        RECT 263.345 66.580 266.140 66.600 ;
        RECT 271.900 66.770 272.430 67.050 ;
        RECT 274.570 66.770 274.740 68.180 ;
        RECT 271.900 66.600 274.740 66.770 ;
        RECT 271.900 66.580 272.410 66.600 ;
        RECT 263.345 65.690 265.825 66.580 ;
        RECT 263.345 64.280 263.515 65.690 ;
        RECT 263.885 65.120 264.925 65.290 ;
        RECT 265.655 64.280 265.825 65.690 ;
        RECT 263.345 64.110 265.825 64.280 ;
      LAYER mcon ;
        RECT 266.310 97.910 266.480 98.080 ;
        RECT 264.455 67.170 264.625 67.340 ;
        RECT 264.815 67.170 264.985 67.340 ;
        RECT 265.930 67.200 266.460 67.730 ;
        RECT 271.580 67.200 272.110 67.730 ;
        RECT 273.055 67.170 273.225 67.340 ;
        RECT 273.415 67.170 273.585 67.340 ;
        RECT 264.140 65.120 264.310 65.290 ;
        RECT 264.500 65.120 264.670 65.290 ;
      LAYER met1 ;
        RECT 266.185 97.955 266.605 98.110 ;
        RECT 268.975 97.955 269.780 98.185 ;
        RECT 266.170 97.580 269.780 97.955 ;
        RECT 268.975 97.300 269.780 97.580 ;
        RECT 264.220 67.200 265.220 67.370 ;
        RECT 265.600 67.200 266.600 68.520 ;
        RECT 264.220 66.970 266.600 67.200 ;
        RECT 265.600 66.130 266.600 66.970 ;
        RECT 271.440 67.200 272.440 68.520 ;
        RECT 272.820 67.200 273.820 67.370 ;
        RECT 271.440 66.970 273.820 67.200 ;
        RECT 271.440 66.130 272.440 66.970 ;
        RECT 265.645 65.540 266.645 66.130 ;
        RECT 263.925 65.320 266.645 65.540 ;
        RECT 263.905 65.275 266.645 65.320 ;
        RECT 263.905 65.090 264.905 65.275 ;
      LAYER via ;
        RECT 269.090 97.455 269.670 98.035 ;
        RECT 265.850 67.365 266.430 68.265 ;
        RECT 271.705 66.340 272.285 66.920 ;
      LAYER met2 ;
        RECT 268.975 98.135 269.780 98.180 ;
        RECT 268.925 97.350 269.830 98.135 ;
        RECT 265.655 67.875 266.645 68.530 ;
        RECT 268.975 67.875 269.780 97.350 ;
        RECT 265.655 67.125 273.000 67.875 ;
        RECT 265.665 67.045 273.000 67.125 ;
        RECT 271.500 66.215 273.000 67.045 ;
        RECT 272.000 63.930 273.000 66.215 ;
      LAYER via2 ;
        RECT 272.200 64.300 272.880 67.820 ;
      LAYER met3 ;
        RECT 272.000 63.930 273.000 67.875 ;
      LAYER via3 ;
        RECT 272.180 64.280 272.900 67.840 ;
      LAYER met4 ;
        RECT 271.670 3.300 273.270 211.800 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 257.010 74.430 257.750 80.460 ;
        RECT 280.290 74.430 281.030 80.460 ;
      LAYER li1 ;
        RECT 205.335 130.980 207.495 131.330 ;
        RECT 252.335 130.980 254.495 131.330 ;
        RECT 283.225 131.200 285.385 131.550 ;
        RECT 205.335 130.150 207.495 130.500 ;
        RECT 252.335 130.150 254.495 130.500 ;
        RECT 257.395 130.060 259.555 130.750 ;
        RECT 278.395 130.060 280.555 130.750 ;
        RECT 283.225 130.370 285.385 130.720 ;
        RECT 330.225 130.370 332.385 130.720 ;
        RECT 205.335 129.320 207.495 129.670 ;
        RECT 252.335 129.320 254.495 129.670 ;
        RECT 257.395 128.890 259.555 129.580 ;
        RECT 278.395 128.890 280.555 129.580 ;
        RECT 283.225 129.540 285.385 129.890 ;
        RECT 330.225 129.540 332.385 129.890 ;
        RECT 205.335 128.490 207.495 128.840 ;
        RECT 252.335 128.490 254.495 128.840 ;
        RECT 283.225 128.710 285.385 129.060 ;
        RECT 330.225 128.710 332.385 129.060 ;
        RECT 205.335 127.660 207.495 128.010 ;
        RECT 252.335 127.660 254.495 128.010 ;
        RECT 257.395 127.720 259.555 128.410 ;
        RECT 278.395 127.720 280.555 128.410 ;
        RECT 283.225 127.880 285.385 128.230 ;
        RECT 330.225 127.880 332.385 128.230 ;
        RECT 205.335 126.830 207.495 127.180 ;
        RECT 252.335 126.830 254.495 127.180 ;
        RECT 257.395 126.550 259.555 127.240 ;
        RECT 278.395 126.550 280.555 127.240 ;
        RECT 283.225 127.050 285.385 127.400 ;
        RECT 330.225 127.050 332.385 127.400 ;
        RECT 205.335 126.000 207.495 126.350 ;
        RECT 252.335 126.000 254.495 126.350 ;
        RECT 283.225 126.220 285.385 126.570 ;
        RECT 330.225 126.220 332.385 126.570 ;
        RECT 205.335 125.170 207.495 125.520 ;
        RECT 252.335 125.170 254.495 125.520 ;
        RECT 257.395 125.380 259.555 126.070 ;
        RECT 278.395 125.380 280.555 126.070 ;
        RECT 283.225 125.390 285.385 125.740 ;
        RECT 330.225 125.390 332.385 125.740 ;
        RECT 205.335 124.340 207.495 124.690 ;
        RECT 252.335 124.340 254.495 124.690 ;
        RECT 257.395 124.210 259.555 124.900 ;
        RECT 278.395 124.210 280.555 124.900 ;
        RECT 283.225 124.560 285.385 124.910 ;
        RECT 330.225 124.560 332.385 124.910 ;
        RECT 205.335 123.510 207.495 123.860 ;
        RECT 252.335 123.510 254.495 123.860 ;
        RECT 283.225 123.730 285.385 124.080 ;
        RECT 330.225 123.730 332.385 124.080 ;
        RECT 257.395 123.040 259.555 123.730 ;
        RECT 278.395 123.040 280.555 123.730 ;
        RECT 205.335 122.680 207.495 123.030 ;
        RECT 252.335 122.680 254.495 123.030 ;
        RECT 283.225 122.900 285.385 123.250 ;
        RECT 330.225 122.900 332.385 123.250 ;
        RECT 205.335 121.850 207.495 122.200 ;
        RECT 252.335 121.850 254.495 122.200 ;
        RECT 257.395 121.870 259.555 122.560 ;
        RECT 278.395 121.870 280.555 122.560 ;
        RECT 283.225 122.070 285.385 122.420 ;
        RECT 330.225 122.070 332.385 122.420 ;
        RECT 205.335 121.020 207.495 121.370 ;
        RECT 252.335 121.020 254.495 121.370 ;
        RECT 257.395 120.700 259.555 121.390 ;
        RECT 278.395 120.700 280.555 121.390 ;
        RECT 283.225 121.240 285.385 121.590 ;
        RECT 330.225 121.240 332.385 121.590 ;
        RECT 205.335 120.190 207.495 120.540 ;
        RECT 252.335 120.190 254.495 120.540 ;
        RECT 283.225 120.410 285.385 120.760 ;
        RECT 330.225 120.410 332.385 120.760 ;
        RECT 205.335 119.360 207.495 119.710 ;
        RECT 252.335 119.360 254.495 119.710 ;
        RECT 257.395 119.530 259.555 120.220 ;
        RECT 278.395 119.530 280.555 120.220 ;
        RECT 283.225 119.580 285.385 119.930 ;
        RECT 330.225 119.580 332.385 119.930 ;
        RECT 205.335 118.530 207.495 118.880 ;
        RECT 252.335 118.530 254.495 118.880 ;
        RECT 257.395 118.360 259.555 119.050 ;
        RECT 278.395 118.360 280.555 119.050 ;
        RECT 283.225 118.750 285.385 119.100 ;
        RECT 330.225 118.750 332.385 119.100 ;
        RECT 205.335 117.700 207.495 118.050 ;
        RECT 252.335 117.700 254.495 118.050 ;
        RECT 283.225 117.920 285.385 118.270 ;
        RECT 330.225 117.920 332.385 118.270 ;
        RECT 205.335 116.870 207.495 117.220 ;
        RECT 252.335 116.870 254.495 117.220 ;
        RECT 257.395 117.190 259.555 117.880 ;
        RECT 278.395 117.190 280.555 117.880 ;
        RECT 283.225 117.090 285.385 117.440 ;
        RECT 330.225 117.090 332.385 117.440 ;
        RECT 205.335 116.040 207.495 116.390 ;
        RECT 252.335 116.040 254.495 116.390 ;
        RECT 257.395 116.020 259.555 116.710 ;
        RECT 278.395 116.020 280.555 116.710 ;
        RECT 283.225 116.260 285.385 116.610 ;
        RECT 330.225 116.260 332.385 116.610 ;
        RECT 205.335 115.210 207.495 115.560 ;
        RECT 252.335 115.210 254.495 115.560 ;
        RECT 257.395 114.850 259.555 115.540 ;
        RECT 278.395 114.850 280.555 115.540 ;
        RECT 283.225 115.430 285.385 115.780 ;
        RECT 330.225 115.430 332.385 115.780 ;
        RECT 205.335 114.380 207.495 114.730 ;
        RECT 252.335 114.380 254.495 114.730 ;
        RECT 283.225 114.600 285.385 114.950 ;
        RECT 330.225 114.600 332.385 114.950 ;
        RECT 205.335 113.550 207.495 113.900 ;
        RECT 252.335 113.550 254.495 113.900 ;
        RECT 257.395 113.680 259.555 114.370 ;
        RECT 278.395 113.680 280.555 114.370 ;
        RECT 283.225 113.770 285.385 114.120 ;
        RECT 330.225 113.770 332.385 114.120 ;
        RECT 205.335 112.720 207.495 113.070 ;
        RECT 252.335 112.720 254.495 113.070 ;
        RECT 257.395 112.510 259.555 113.200 ;
        RECT 278.395 112.510 280.555 113.200 ;
        RECT 283.225 112.940 285.385 113.290 ;
        RECT 330.225 112.940 332.385 113.290 ;
        RECT 205.335 111.890 207.495 112.240 ;
        RECT 252.335 111.890 254.495 112.240 ;
        RECT 283.225 112.110 285.385 112.460 ;
        RECT 330.225 112.110 332.385 112.460 ;
        RECT 205.335 111.060 207.495 111.410 ;
        RECT 252.335 111.060 254.495 111.410 ;
        RECT 257.395 111.340 259.555 112.030 ;
        RECT 278.395 111.340 280.555 112.030 ;
        RECT 283.225 111.280 285.385 111.630 ;
        RECT 330.225 111.280 332.385 111.630 ;
        RECT 205.335 110.230 207.495 110.580 ;
        RECT 252.335 110.230 254.495 110.580 ;
        RECT 257.395 110.170 259.555 110.860 ;
        RECT 278.395 110.170 280.555 110.860 ;
        RECT 283.225 110.450 285.385 110.800 ;
        RECT 330.225 110.450 332.385 110.800 ;
        RECT 205.335 109.400 207.495 109.750 ;
        RECT 252.335 109.400 254.495 109.750 ;
        RECT 257.395 109.000 259.555 109.690 ;
        RECT 278.395 109.000 280.555 109.690 ;
        RECT 283.225 109.620 285.385 109.970 ;
        RECT 330.225 109.620 332.385 109.970 ;
        RECT 205.335 108.570 207.495 108.920 ;
        RECT 252.335 108.570 254.495 108.920 ;
        RECT 283.225 108.790 285.385 109.140 ;
        RECT 330.225 108.790 332.385 109.140 ;
        RECT 205.335 107.740 207.495 108.090 ;
        RECT 252.335 107.740 254.495 108.090 ;
        RECT 257.395 107.830 259.555 108.520 ;
        RECT 278.395 107.830 280.555 108.520 ;
        RECT 283.225 107.960 285.385 108.310 ;
        RECT 330.225 107.960 332.385 108.310 ;
        RECT 205.335 106.910 207.495 107.260 ;
        RECT 252.335 106.910 254.495 107.260 ;
        RECT 257.395 106.660 259.555 107.350 ;
        RECT 278.395 106.660 280.555 107.350 ;
        RECT 283.225 107.130 285.385 107.480 ;
        RECT 330.225 107.130 332.385 107.480 ;
        RECT 205.335 106.080 207.495 106.430 ;
        RECT 252.335 106.080 254.495 106.430 ;
        RECT 283.225 106.300 285.385 106.650 ;
        RECT 330.225 106.300 332.385 106.650 ;
        RECT 205.335 105.250 207.495 105.600 ;
        RECT 252.335 105.250 254.495 105.600 ;
        RECT 257.395 105.490 259.555 106.180 ;
        RECT 278.395 105.490 280.555 106.180 ;
        RECT 283.225 105.470 285.385 105.820 ;
        RECT 330.225 105.470 332.385 105.820 ;
        RECT 205.335 104.420 207.495 104.770 ;
        RECT 252.335 104.420 254.495 104.770 ;
        RECT 257.395 104.320 259.555 105.010 ;
        RECT 278.395 104.320 280.555 105.010 ;
        RECT 283.225 104.640 285.385 104.990 ;
        RECT 330.225 104.640 332.385 104.990 ;
        RECT 205.335 103.590 207.495 103.940 ;
        RECT 252.335 103.590 254.495 103.940 ;
        RECT 257.395 103.150 259.555 103.840 ;
        RECT 278.395 103.150 280.555 103.840 ;
        RECT 283.225 103.810 285.385 104.160 ;
        RECT 330.225 103.810 332.385 104.160 ;
        RECT 205.335 102.760 207.495 103.110 ;
        RECT 252.335 102.760 254.495 103.110 ;
        RECT 283.225 102.980 285.385 103.330 ;
        RECT 330.225 102.980 332.385 103.330 ;
        RECT 205.335 101.930 207.495 102.280 ;
        RECT 252.335 101.930 254.495 102.280 ;
        RECT 283.225 102.150 285.385 102.500 ;
        RECT 330.225 102.150 332.385 102.500 ;
        RECT 205.335 101.100 207.495 101.450 ;
        RECT 252.335 101.100 254.495 101.450 ;
        RECT 283.225 101.320 285.385 101.670 ;
        RECT 330.225 101.320 332.385 101.670 ;
        RECT 205.335 100.270 207.495 100.620 ;
        RECT 252.335 100.270 254.495 100.620 ;
        RECT 283.225 100.490 285.385 100.840 ;
        RECT 330.225 100.490 332.385 100.840 ;
        RECT 205.335 99.440 207.495 99.790 ;
        RECT 252.335 99.440 254.495 99.790 ;
        RECT 283.225 99.660 285.385 100.010 ;
        RECT 330.225 99.660 332.385 100.010 ;
        RECT 270.455 99.180 270.915 99.350 ;
        RECT 273.145 99.180 273.605 99.350 ;
        RECT 205.335 98.610 207.495 98.960 ;
        RECT 252.335 98.610 254.495 98.960 ;
        RECT 266.165 98.700 266.625 98.870 ;
        RECT 266.840 98.140 267.010 98.640 ;
        RECT 270.115 98.620 270.285 99.120 ;
        RECT 273.775 98.620 273.945 99.120 ;
        RECT 283.225 98.830 285.385 99.180 ;
        RECT 330.225 98.830 332.385 99.180 ;
        RECT 270.455 98.390 270.915 98.560 ;
        RECT 205.335 97.780 207.495 98.130 ;
        RECT 252.335 97.780 254.495 98.130 ;
        RECT 283.225 98.000 285.385 98.350 ;
        RECT 330.225 98.000 332.385 98.350 ;
        RECT 205.335 96.950 207.495 97.300 ;
        RECT 252.335 96.950 254.495 97.300 ;
        RECT 283.225 97.170 285.385 97.520 ;
        RECT 330.225 97.170 332.385 97.520 ;
        RECT 205.335 96.120 207.495 96.470 ;
        RECT 252.335 96.120 254.495 96.470 ;
        RECT 270.455 96.400 270.915 96.570 ;
        RECT 273.145 96.400 273.605 96.570 ;
        RECT 283.225 96.340 285.385 96.690 ;
        RECT 330.225 96.340 332.385 96.690 ;
        RECT 270.115 95.840 270.285 96.340 ;
        RECT 273.775 95.840 273.945 96.340 ;
        RECT 205.335 95.290 207.495 95.640 ;
        RECT 252.335 95.290 254.495 95.640 ;
        RECT 266.165 95.620 266.625 95.790 ;
        RECT 270.455 95.610 270.915 95.780 ;
        RECT 262.750 95.060 262.920 95.560 ;
        RECT 266.840 95.060 267.010 95.560 ;
        RECT 283.225 95.510 285.385 95.860 ;
        RECT 330.225 95.510 332.385 95.860 ;
        RECT 263.135 94.830 263.595 95.000 ;
        RECT 266.165 94.830 266.625 95.000 ;
        RECT 205.335 94.460 207.495 94.810 ;
        RECT 252.335 94.460 254.495 94.810 ;
        RECT 283.225 94.680 285.385 95.030 ;
        RECT 330.225 94.680 332.385 95.030 ;
        RECT 205.335 93.630 207.495 93.980 ;
        RECT 252.335 93.630 254.495 93.980 ;
        RECT 283.225 93.850 285.385 94.200 ;
        RECT 330.225 93.850 332.385 94.200 ;
        RECT 270.455 93.620 270.915 93.790 ;
        RECT 273.145 93.620 273.605 93.790 ;
        RECT 276.775 93.610 277.235 93.780 ;
        RECT 205.335 92.800 207.495 93.150 ;
        RECT 252.335 92.800 254.495 93.150 ;
        RECT 270.115 93.060 270.285 93.560 ;
        RECT 273.775 93.060 273.945 93.560 ;
        RECT 277.405 93.050 277.575 93.550 ;
        RECT 283.225 93.020 285.385 93.370 ;
        RECT 330.225 93.020 332.385 93.370 ;
        RECT 270.455 92.830 270.915 93.000 ;
        RECT 266.165 92.540 266.625 92.710 ;
        RECT 205.335 91.970 207.495 92.320 ;
        RECT 252.335 91.970 254.495 92.320 ;
        RECT 262.750 91.980 262.920 92.480 ;
        RECT 266.840 91.980 267.010 92.480 ;
        RECT 283.225 92.190 285.385 92.540 ;
        RECT 330.225 92.190 332.385 92.540 ;
        RECT 263.135 91.750 263.595 91.920 ;
        RECT 266.165 91.750 266.625 91.920 ;
        RECT 205.335 91.140 207.495 91.490 ;
        RECT 252.335 91.140 254.495 91.490 ;
        RECT 283.225 91.360 285.385 91.710 ;
        RECT 330.225 91.360 332.385 91.710 ;
        RECT 270.455 90.840 270.915 91.010 ;
        RECT 273.145 90.840 273.605 91.010 ;
        RECT 205.335 90.310 207.495 90.660 ;
        RECT 252.335 90.310 254.495 90.660 ;
        RECT 273.775 90.280 273.945 90.780 ;
        RECT 277.405 90.270 277.575 90.770 ;
        RECT 283.225 90.530 285.385 90.880 ;
        RECT 330.225 90.530 332.385 90.880 ;
        RECT 270.455 90.050 270.915 90.220 ;
        RECT 205.335 89.480 207.495 89.830 ;
        RECT 252.335 89.480 254.495 89.830 ;
        RECT 283.225 89.700 285.385 90.050 ;
        RECT 330.225 89.700 332.385 90.050 ;
        RECT 266.165 89.460 266.625 89.630 ;
        RECT 205.335 88.650 207.495 89.000 ;
        RECT 252.335 88.650 254.495 89.000 ;
        RECT 262.750 88.900 262.920 89.400 ;
        RECT 283.225 88.870 285.385 89.220 ;
        RECT 330.225 88.870 332.385 89.220 ;
        RECT 263.135 88.670 263.595 88.840 ;
        RECT 266.165 88.670 266.625 88.840 ;
        RECT 205.335 87.820 207.495 88.170 ;
        RECT 252.335 87.820 254.495 88.170 ;
        RECT 270.455 88.060 270.915 88.230 ;
        RECT 273.145 88.060 273.605 88.230 ;
        RECT 276.775 88.050 277.235 88.220 ;
        RECT 283.225 88.040 285.385 88.390 ;
        RECT 330.225 88.040 332.385 88.390 ;
        RECT 270.115 87.500 270.285 88.000 ;
        RECT 273.775 87.500 273.945 88.000 ;
        RECT 277.405 87.490 277.575 87.990 ;
        RECT 205.335 86.990 207.495 87.340 ;
        RECT 252.335 86.990 254.495 87.340 ;
        RECT 270.455 87.270 270.915 87.440 ;
        RECT 283.225 87.210 285.385 87.560 ;
        RECT 330.225 87.210 332.385 87.560 ;
        RECT 205.335 86.160 207.495 86.510 ;
        RECT 252.335 86.160 254.495 86.510 ;
        RECT 263.135 86.380 263.595 86.550 ;
        RECT 266.165 86.380 266.625 86.550 ;
        RECT 283.225 86.380 285.385 86.730 ;
        RECT 330.225 86.380 332.385 86.730 ;
        RECT 262.750 85.820 262.920 86.320 ;
        RECT 266.840 85.820 267.010 86.320 ;
        RECT 205.335 85.330 207.495 85.680 ;
        RECT 252.335 85.330 254.495 85.680 ;
        RECT 283.225 85.550 285.385 85.900 ;
        RECT 330.225 85.550 332.385 85.900 ;
        RECT 270.455 85.280 270.915 85.450 ;
        RECT 273.145 85.280 273.605 85.450 ;
        RECT 276.775 85.270 277.235 85.440 ;
        RECT 252.335 84.500 254.495 84.850 ;
        RECT 270.115 84.720 270.285 85.220 ;
        RECT 273.775 84.720 273.945 85.220 ;
        RECT 277.405 84.710 277.575 85.210 ;
        RECT 283.225 84.720 285.385 85.070 ;
        RECT 330.225 84.720 332.385 85.070 ;
        RECT 270.455 84.490 270.915 84.660 ;
        RECT 276.775 84.480 277.235 84.650 ;
        RECT 283.225 83.890 285.385 84.240 ;
        RECT 330.225 83.890 332.385 84.240 ;
        RECT 283.225 83.060 285.385 83.410 ;
        RECT 330.225 83.060 332.385 83.410 ;
        RECT 283.225 82.230 285.385 82.580 ;
        RECT 330.225 82.230 332.385 82.580 ;
        RECT 205.385 81.500 207.545 81.850 ;
        RECT 252.385 81.500 254.545 81.850 ;
        RECT 283.225 81.400 285.385 81.750 ;
        RECT 330.225 81.400 332.385 81.750 ;
        RECT 205.385 80.670 207.545 81.020 ;
        RECT 252.385 80.670 254.545 81.020 ;
        RECT 283.225 80.570 285.385 80.920 ;
        RECT 330.225 80.570 332.385 80.920 ;
        RECT 205.385 79.840 207.545 80.190 ;
        RECT 252.385 79.840 254.545 80.190 ;
        RECT 205.385 79.010 207.545 79.360 ;
        RECT 252.385 79.010 254.545 79.360 ;
        RECT 205.385 78.180 207.545 78.530 ;
        RECT 252.385 78.180 254.545 78.530 ;
        RECT 205.385 77.350 207.545 77.700 ;
        RECT 252.385 77.350 254.545 77.700 ;
        RECT 205.385 76.520 207.545 76.870 ;
        RECT 252.385 76.520 254.545 76.870 ;
        RECT 205.385 75.690 207.545 76.040 ;
        RECT 252.385 75.690 254.545 76.040 ;
        RECT 205.385 74.860 207.545 75.210 ;
        RECT 252.385 74.860 254.545 75.210 ;
        RECT 257.140 74.600 257.620 80.290 ;
        RECT 263.185 79.100 263.645 79.270 ;
        RECT 266.535 79.100 266.995 79.270 ;
        RECT 271.045 79.100 271.505 79.270 ;
        RECT 274.395 79.100 274.855 79.270 ;
        RECT 259.350 78.530 259.520 79.030 ;
        RECT 260.320 78.530 260.490 79.030 ;
        RECT 262.800 78.540 262.970 79.040 ;
        RECT 263.860 78.540 264.030 79.040 ;
        RECT 266.150 78.540 266.320 79.040 ;
        RECT 267.210 78.540 267.380 79.040 ;
        RECT 270.660 78.540 270.830 79.040 ;
        RECT 271.720 78.540 271.890 79.040 ;
        RECT 274.010 78.540 274.180 79.040 ;
        RECT 275.070 78.540 275.240 79.040 ;
        RECT 277.550 78.530 277.720 79.030 ;
        RECT 278.520 78.530 278.690 79.030 ;
        RECT 259.690 78.300 260.150 78.470 ;
        RECT 263.185 78.310 263.645 78.480 ;
        RECT 274.395 78.310 274.855 78.480 ;
        RECT 277.890 78.300 278.350 78.470 ;
        RECT 259.680 76.060 260.140 76.230 ;
        RECT 263.195 76.050 263.655 76.220 ;
        RECT 274.385 76.050 274.845 76.220 ;
        RECT 277.900 76.060 278.360 76.230 ;
        RECT 262.810 75.490 262.980 75.990 ;
        RECT 263.870 75.490 264.040 75.990 ;
        RECT 266.150 75.460 266.320 75.960 ;
        RECT 267.210 75.460 267.380 75.960 ;
        RECT 270.660 75.460 270.830 75.960 ;
        RECT 271.720 75.460 271.890 75.960 ;
        RECT 274.000 75.490 274.170 75.990 ;
        RECT 275.060 75.490 275.230 75.990 ;
        RECT 263.195 75.260 263.655 75.430 ;
        RECT 266.535 75.230 266.995 75.400 ;
        RECT 271.045 75.230 271.505 75.400 ;
        RECT 274.385 75.260 274.845 75.430 ;
        RECT 280.420 74.600 280.900 80.290 ;
        RECT 283.225 79.740 285.385 80.090 ;
        RECT 330.225 79.740 332.385 80.090 ;
        RECT 283.225 78.910 285.385 79.260 ;
        RECT 330.225 78.910 332.385 79.260 ;
        RECT 283.225 78.080 285.385 78.430 ;
        RECT 330.225 78.080 332.385 78.430 ;
        RECT 283.225 77.250 285.385 77.600 ;
        RECT 330.225 77.250 332.385 77.600 ;
        RECT 283.225 76.420 285.385 76.770 ;
        RECT 330.225 76.420 332.385 76.770 ;
        RECT 283.225 75.590 285.385 75.940 ;
        RECT 330.225 75.590 332.385 75.940 ;
        RECT 283.225 74.760 285.385 75.110 ;
        RECT 330.225 74.760 332.385 75.110 ;
        RECT 205.385 74.030 207.545 74.380 ;
        RECT 252.385 74.030 254.545 74.380 ;
        RECT 283.225 73.930 285.385 74.280 ;
        RECT 330.225 73.930 332.385 74.280 ;
        RECT 205.385 73.200 207.545 73.550 ;
        RECT 252.385 73.200 254.545 73.550 ;
        RECT 283.225 73.100 285.385 73.450 ;
        RECT 330.225 73.100 332.385 73.450 ;
        RECT 205.385 72.370 207.545 72.720 ;
        RECT 252.385 72.370 254.545 72.720 ;
        RECT 283.225 72.270 285.385 72.620 ;
        RECT 330.225 72.270 332.385 72.620 ;
        RECT 205.385 71.540 207.545 71.890 ;
        RECT 252.385 71.540 254.545 71.890 ;
        RECT 283.225 71.440 285.385 71.790 ;
        RECT 330.225 71.440 332.385 71.790 ;
        RECT 205.385 70.710 207.545 71.060 ;
        RECT 252.385 70.710 254.545 71.060 ;
        RECT 274.025 70.320 276.185 71.010 ;
        RECT 283.225 70.610 285.385 70.960 ;
        RECT 330.225 70.610 332.385 70.960 ;
        RECT 205.385 69.880 207.545 70.230 ;
        RECT 252.385 69.880 254.545 70.230 ;
        RECT 283.225 69.780 285.385 70.130 ;
        RECT 330.225 69.780 332.385 70.130 ;
        RECT 205.385 69.050 207.545 69.400 ;
        RECT 252.385 69.050 254.545 69.400 ;
        RECT 283.225 68.950 285.385 69.300 ;
        RECT 330.225 68.950 332.385 69.300 ;
        RECT 205.385 68.220 207.545 68.570 ;
        RECT 252.385 68.220 254.545 68.570 ;
        RECT 283.225 68.120 285.385 68.470 ;
        RECT 330.225 68.120 332.385 68.470 ;
        RECT 205.385 67.390 207.545 67.740 ;
        RECT 252.385 67.390 254.545 67.740 ;
        RECT 261.010 67.610 262.050 67.780 ;
        RECT 264.200 67.610 265.240 67.780 ;
        RECT 272.800 67.610 273.840 67.780 ;
        RECT 275.990 67.610 277.030 67.780 ;
        RECT 283.225 67.290 285.385 67.640 ;
        RECT 330.225 67.290 332.385 67.640 ;
        RECT 252.385 66.560 254.545 66.910 ;
        RECT 267.885 66.885 268.055 67.215 ;
        RECT 268.225 66.745 268.765 66.915 ;
        RECT 283.225 66.460 285.385 66.810 ;
        RECT 330.225 66.460 332.385 66.810 ;
        RECT 263.885 64.680 264.925 64.850 ;
        RECT 265.140 64.820 265.310 65.150 ;
        RECT 268.225 65.120 268.765 65.290 ;
        RECT 268.225 64.680 268.765 64.850 ;
        RECT 270.175 64.820 270.345 65.150 ;
        RECT 270.515 64.680 270.975 64.850 ;
      LAYER mcon ;
        RECT 205.435 131.070 205.605 131.240 ;
        RECT 205.795 131.070 205.965 131.240 ;
        RECT 206.155 131.070 206.325 131.240 ;
        RECT 206.515 131.070 206.685 131.240 ;
        RECT 206.875 131.070 207.045 131.240 ;
        RECT 207.235 131.070 207.405 131.240 ;
        RECT 252.430 131.070 252.600 131.240 ;
        RECT 252.790 131.070 252.960 131.240 ;
        RECT 253.150 131.070 253.320 131.240 ;
        RECT 253.510 131.070 253.680 131.240 ;
        RECT 253.870 131.070 254.040 131.240 ;
        RECT 254.230 131.070 254.400 131.240 ;
        RECT 283.325 131.290 283.495 131.460 ;
        RECT 283.685 131.290 283.855 131.460 ;
        RECT 284.045 131.290 284.215 131.460 ;
        RECT 284.405 131.290 284.575 131.460 ;
        RECT 284.765 131.290 284.935 131.460 ;
        RECT 285.125 131.290 285.295 131.460 ;
        RECT 205.435 130.240 205.605 130.410 ;
        RECT 205.795 130.240 205.965 130.410 ;
        RECT 206.155 130.240 206.325 130.410 ;
        RECT 206.515 130.240 206.685 130.410 ;
        RECT 206.875 130.240 207.045 130.410 ;
        RECT 207.235 130.240 207.405 130.410 ;
        RECT 252.430 130.240 252.600 130.410 ;
        RECT 252.790 130.240 252.960 130.410 ;
        RECT 253.150 130.240 253.320 130.410 ;
        RECT 253.510 130.240 253.680 130.410 ;
        RECT 253.870 130.240 254.040 130.410 ;
        RECT 254.230 130.240 254.400 130.410 ;
        RECT 257.495 130.140 259.465 130.670 ;
        RECT 278.490 130.140 280.460 130.670 ;
        RECT 283.325 130.460 283.495 130.630 ;
        RECT 283.685 130.460 283.855 130.630 ;
        RECT 284.045 130.460 284.215 130.630 ;
        RECT 284.405 130.460 284.575 130.630 ;
        RECT 284.765 130.460 284.935 130.630 ;
        RECT 285.125 130.460 285.295 130.630 ;
        RECT 330.320 130.460 330.490 130.630 ;
        RECT 330.680 130.460 330.850 130.630 ;
        RECT 331.040 130.460 331.210 130.630 ;
        RECT 331.400 130.460 331.570 130.630 ;
        RECT 331.760 130.460 331.930 130.630 ;
        RECT 332.120 130.460 332.290 130.630 ;
        RECT 205.435 129.410 205.605 129.580 ;
        RECT 205.795 129.410 205.965 129.580 ;
        RECT 206.155 129.410 206.325 129.580 ;
        RECT 206.515 129.410 206.685 129.580 ;
        RECT 206.875 129.410 207.045 129.580 ;
        RECT 207.235 129.410 207.405 129.580 ;
        RECT 283.325 129.630 283.495 129.800 ;
        RECT 283.685 129.630 283.855 129.800 ;
        RECT 284.045 129.630 284.215 129.800 ;
        RECT 284.405 129.630 284.575 129.800 ;
        RECT 284.765 129.630 284.935 129.800 ;
        RECT 285.125 129.630 285.295 129.800 ;
        RECT 252.430 129.410 252.600 129.580 ;
        RECT 252.790 129.410 252.960 129.580 ;
        RECT 253.150 129.410 253.320 129.580 ;
        RECT 253.510 129.410 253.680 129.580 ;
        RECT 253.870 129.410 254.040 129.580 ;
        RECT 254.230 129.410 254.400 129.580 ;
        RECT 257.495 128.970 259.465 129.500 ;
        RECT 330.320 129.630 330.490 129.800 ;
        RECT 330.680 129.630 330.850 129.800 ;
        RECT 331.040 129.630 331.210 129.800 ;
        RECT 331.400 129.630 331.570 129.800 ;
        RECT 331.760 129.630 331.930 129.800 ;
        RECT 332.120 129.630 332.290 129.800 ;
        RECT 278.490 128.970 280.460 129.500 ;
        RECT 205.435 128.580 205.605 128.750 ;
        RECT 205.795 128.580 205.965 128.750 ;
        RECT 206.155 128.580 206.325 128.750 ;
        RECT 206.515 128.580 206.685 128.750 ;
        RECT 206.875 128.580 207.045 128.750 ;
        RECT 207.235 128.580 207.405 128.750 ;
        RECT 252.430 128.580 252.600 128.750 ;
        RECT 252.790 128.580 252.960 128.750 ;
        RECT 253.150 128.580 253.320 128.750 ;
        RECT 253.510 128.580 253.680 128.750 ;
        RECT 253.870 128.580 254.040 128.750 ;
        RECT 254.230 128.580 254.400 128.750 ;
        RECT 283.325 128.800 283.495 128.970 ;
        RECT 283.685 128.800 283.855 128.970 ;
        RECT 284.045 128.800 284.215 128.970 ;
        RECT 284.405 128.800 284.575 128.970 ;
        RECT 284.765 128.800 284.935 128.970 ;
        RECT 285.125 128.800 285.295 128.970 ;
        RECT 330.320 128.800 330.490 128.970 ;
        RECT 330.680 128.800 330.850 128.970 ;
        RECT 331.040 128.800 331.210 128.970 ;
        RECT 331.400 128.800 331.570 128.970 ;
        RECT 331.760 128.800 331.930 128.970 ;
        RECT 332.120 128.800 332.290 128.970 ;
        RECT 205.435 127.750 205.605 127.920 ;
        RECT 205.795 127.750 205.965 127.920 ;
        RECT 206.155 127.750 206.325 127.920 ;
        RECT 206.515 127.750 206.685 127.920 ;
        RECT 206.875 127.750 207.045 127.920 ;
        RECT 207.235 127.750 207.405 127.920 ;
        RECT 252.430 127.750 252.600 127.920 ;
        RECT 252.790 127.750 252.960 127.920 ;
        RECT 253.150 127.750 253.320 127.920 ;
        RECT 253.510 127.750 253.680 127.920 ;
        RECT 253.870 127.750 254.040 127.920 ;
        RECT 254.230 127.750 254.400 127.920 ;
        RECT 257.495 127.800 259.465 128.330 ;
        RECT 278.490 127.800 280.460 128.330 ;
        RECT 283.325 127.970 283.495 128.140 ;
        RECT 283.685 127.970 283.855 128.140 ;
        RECT 284.045 127.970 284.215 128.140 ;
        RECT 284.405 127.970 284.575 128.140 ;
        RECT 284.765 127.970 284.935 128.140 ;
        RECT 285.125 127.970 285.295 128.140 ;
        RECT 330.320 127.970 330.490 128.140 ;
        RECT 330.680 127.970 330.850 128.140 ;
        RECT 331.040 127.970 331.210 128.140 ;
        RECT 331.400 127.970 331.570 128.140 ;
        RECT 331.760 127.970 331.930 128.140 ;
        RECT 332.120 127.970 332.290 128.140 ;
        RECT 205.435 126.920 205.605 127.090 ;
        RECT 205.795 126.920 205.965 127.090 ;
        RECT 206.155 126.920 206.325 127.090 ;
        RECT 206.515 126.920 206.685 127.090 ;
        RECT 206.875 126.920 207.045 127.090 ;
        RECT 207.235 126.920 207.405 127.090 ;
        RECT 252.430 126.920 252.600 127.090 ;
        RECT 252.790 126.920 252.960 127.090 ;
        RECT 253.150 126.920 253.320 127.090 ;
        RECT 253.510 126.920 253.680 127.090 ;
        RECT 253.870 126.920 254.040 127.090 ;
        RECT 254.230 126.920 254.400 127.090 ;
        RECT 257.495 126.630 259.465 127.160 ;
        RECT 278.490 126.630 280.460 127.160 ;
        RECT 283.325 127.140 283.495 127.310 ;
        RECT 283.685 127.140 283.855 127.310 ;
        RECT 284.045 127.140 284.215 127.310 ;
        RECT 284.405 127.140 284.575 127.310 ;
        RECT 284.765 127.140 284.935 127.310 ;
        RECT 285.125 127.140 285.295 127.310 ;
        RECT 330.320 127.140 330.490 127.310 ;
        RECT 330.680 127.140 330.850 127.310 ;
        RECT 331.040 127.140 331.210 127.310 ;
        RECT 331.400 127.140 331.570 127.310 ;
        RECT 331.760 127.140 331.930 127.310 ;
        RECT 332.120 127.140 332.290 127.310 ;
        RECT 205.435 126.090 205.605 126.260 ;
        RECT 205.795 126.090 205.965 126.260 ;
        RECT 206.155 126.090 206.325 126.260 ;
        RECT 206.515 126.090 206.685 126.260 ;
        RECT 206.875 126.090 207.045 126.260 ;
        RECT 207.235 126.090 207.405 126.260 ;
        RECT 252.430 126.090 252.600 126.260 ;
        RECT 252.790 126.090 252.960 126.260 ;
        RECT 253.150 126.090 253.320 126.260 ;
        RECT 253.510 126.090 253.680 126.260 ;
        RECT 253.870 126.090 254.040 126.260 ;
        RECT 254.230 126.090 254.400 126.260 ;
        RECT 283.325 126.310 283.495 126.480 ;
        RECT 283.685 126.310 283.855 126.480 ;
        RECT 284.045 126.310 284.215 126.480 ;
        RECT 284.405 126.310 284.575 126.480 ;
        RECT 284.765 126.310 284.935 126.480 ;
        RECT 285.125 126.310 285.295 126.480 ;
        RECT 330.320 126.310 330.490 126.480 ;
        RECT 330.680 126.310 330.850 126.480 ;
        RECT 331.040 126.310 331.210 126.480 ;
        RECT 331.400 126.310 331.570 126.480 ;
        RECT 331.760 126.310 331.930 126.480 ;
        RECT 332.120 126.310 332.290 126.480 ;
        RECT 205.435 125.260 205.605 125.430 ;
        RECT 205.795 125.260 205.965 125.430 ;
        RECT 206.155 125.260 206.325 125.430 ;
        RECT 206.515 125.260 206.685 125.430 ;
        RECT 206.875 125.260 207.045 125.430 ;
        RECT 207.235 125.260 207.405 125.430 ;
        RECT 252.430 125.260 252.600 125.430 ;
        RECT 252.790 125.260 252.960 125.430 ;
        RECT 253.150 125.260 253.320 125.430 ;
        RECT 253.510 125.260 253.680 125.430 ;
        RECT 253.870 125.260 254.040 125.430 ;
        RECT 254.230 125.260 254.400 125.430 ;
        RECT 257.495 125.460 259.465 125.990 ;
        RECT 278.490 125.460 280.460 125.990 ;
        RECT 283.325 125.480 283.495 125.650 ;
        RECT 283.685 125.480 283.855 125.650 ;
        RECT 284.045 125.480 284.215 125.650 ;
        RECT 284.405 125.480 284.575 125.650 ;
        RECT 284.765 125.480 284.935 125.650 ;
        RECT 285.125 125.480 285.295 125.650 ;
        RECT 330.320 125.480 330.490 125.650 ;
        RECT 330.680 125.480 330.850 125.650 ;
        RECT 331.040 125.480 331.210 125.650 ;
        RECT 331.400 125.480 331.570 125.650 ;
        RECT 331.760 125.480 331.930 125.650 ;
        RECT 332.120 125.480 332.290 125.650 ;
        RECT 205.435 124.430 205.605 124.600 ;
        RECT 205.795 124.430 205.965 124.600 ;
        RECT 206.155 124.430 206.325 124.600 ;
        RECT 206.515 124.430 206.685 124.600 ;
        RECT 206.875 124.430 207.045 124.600 ;
        RECT 207.235 124.430 207.405 124.600 ;
        RECT 252.430 124.430 252.600 124.600 ;
        RECT 252.790 124.430 252.960 124.600 ;
        RECT 253.150 124.430 253.320 124.600 ;
        RECT 253.510 124.430 253.680 124.600 ;
        RECT 253.870 124.430 254.040 124.600 ;
        RECT 254.230 124.430 254.400 124.600 ;
        RECT 257.495 124.290 259.465 124.820 ;
        RECT 278.490 124.290 280.460 124.820 ;
        RECT 283.325 124.650 283.495 124.820 ;
        RECT 283.685 124.650 283.855 124.820 ;
        RECT 284.045 124.650 284.215 124.820 ;
        RECT 284.405 124.650 284.575 124.820 ;
        RECT 284.765 124.650 284.935 124.820 ;
        RECT 285.125 124.650 285.295 124.820 ;
        RECT 330.320 124.650 330.490 124.820 ;
        RECT 330.680 124.650 330.850 124.820 ;
        RECT 331.040 124.650 331.210 124.820 ;
        RECT 331.400 124.650 331.570 124.820 ;
        RECT 331.760 124.650 331.930 124.820 ;
        RECT 332.120 124.650 332.290 124.820 ;
        RECT 205.435 123.600 205.605 123.770 ;
        RECT 205.795 123.600 205.965 123.770 ;
        RECT 206.155 123.600 206.325 123.770 ;
        RECT 206.515 123.600 206.685 123.770 ;
        RECT 206.875 123.600 207.045 123.770 ;
        RECT 207.235 123.600 207.405 123.770 ;
        RECT 252.430 123.600 252.600 123.770 ;
        RECT 252.790 123.600 252.960 123.770 ;
        RECT 253.150 123.600 253.320 123.770 ;
        RECT 253.510 123.600 253.680 123.770 ;
        RECT 253.870 123.600 254.040 123.770 ;
        RECT 254.230 123.600 254.400 123.770 ;
        RECT 283.325 123.820 283.495 123.990 ;
        RECT 283.685 123.820 283.855 123.990 ;
        RECT 284.045 123.820 284.215 123.990 ;
        RECT 284.405 123.820 284.575 123.990 ;
        RECT 284.765 123.820 284.935 123.990 ;
        RECT 285.125 123.820 285.295 123.990 ;
        RECT 330.320 123.820 330.490 123.990 ;
        RECT 330.680 123.820 330.850 123.990 ;
        RECT 331.040 123.820 331.210 123.990 ;
        RECT 331.400 123.820 331.570 123.990 ;
        RECT 331.760 123.820 331.930 123.990 ;
        RECT 332.120 123.820 332.290 123.990 ;
        RECT 257.495 123.120 259.465 123.650 ;
        RECT 278.490 123.120 280.460 123.650 ;
        RECT 205.435 122.770 205.605 122.940 ;
        RECT 205.795 122.770 205.965 122.940 ;
        RECT 206.155 122.770 206.325 122.940 ;
        RECT 206.515 122.770 206.685 122.940 ;
        RECT 206.875 122.770 207.045 122.940 ;
        RECT 207.235 122.770 207.405 122.940 ;
        RECT 252.430 122.770 252.600 122.940 ;
        RECT 252.790 122.770 252.960 122.940 ;
        RECT 253.150 122.770 253.320 122.940 ;
        RECT 253.510 122.770 253.680 122.940 ;
        RECT 253.870 122.770 254.040 122.940 ;
        RECT 254.230 122.770 254.400 122.940 ;
        RECT 283.325 122.990 283.495 123.160 ;
        RECT 283.685 122.990 283.855 123.160 ;
        RECT 284.045 122.990 284.215 123.160 ;
        RECT 284.405 122.990 284.575 123.160 ;
        RECT 284.765 122.990 284.935 123.160 ;
        RECT 285.125 122.990 285.295 123.160 ;
        RECT 330.320 122.990 330.490 123.160 ;
        RECT 330.680 122.990 330.850 123.160 ;
        RECT 331.040 122.990 331.210 123.160 ;
        RECT 331.400 122.990 331.570 123.160 ;
        RECT 331.760 122.990 331.930 123.160 ;
        RECT 332.120 122.990 332.290 123.160 ;
        RECT 205.435 121.940 205.605 122.110 ;
        RECT 205.795 121.940 205.965 122.110 ;
        RECT 206.155 121.940 206.325 122.110 ;
        RECT 206.515 121.940 206.685 122.110 ;
        RECT 206.875 121.940 207.045 122.110 ;
        RECT 207.235 121.940 207.405 122.110 ;
        RECT 252.430 121.940 252.600 122.110 ;
        RECT 252.790 121.940 252.960 122.110 ;
        RECT 253.150 121.940 253.320 122.110 ;
        RECT 253.510 121.940 253.680 122.110 ;
        RECT 253.870 121.940 254.040 122.110 ;
        RECT 254.230 121.940 254.400 122.110 ;
        RECT 257.495 121.950 259.465 122.480 ;
        RECT 278.490 121.950 280.460 122.480 ;
        RECT 283.325 122.160 283.495 122.330 ;
        RECT 283.685 122.160 283.855 122.330 ;
        RECT 284.045 122.160 284.215 122.330 ;
        RECT 284.405 122.160 284.575 122.330 ;
        RECT 284.765 122.160 284.935 122.330 ;
        RECT 285.125 122.160 285.295 122.330 ;
        RECT 330.320 122.160 330.490 122.330 ;
        RECT 330.680 122.160 330.850 122.330 ;
        RECT 331.040 122.160 331.210 122.330 ;
        RECT 331.400 122.160 331.570 122.330 ;
        RECT 331.760 122.160 331.930 122.330 ;
        RECT 332.120 122.160 332.290 122.330 ;
        RECT 205.435 121.110 205.605 121.280 ;
        RECT 205.795 121.110 205.965 121.280 ;
        RECT 206.155 121.110 206.325 121.280 ;
        RECT 206.515 121.110 206.685 121.280 ;
        RECT 206.875 121.110 207.045 121.280 ;
        RECT 207.235 121.110 207.405 121.280 ;
        RECT 252.430 121.110 252.600 121.280 ;
        RECT 252.790 121.110 252.960 121.280 ;
        RECT 253.150 121.110 253.320 121.280 ;
        RECT 253.510 121.110 253.680 121.280 ;
        RECT 253.870 121.110 254.040 121.280 ;
        RECT 254.230 121.110 254.400 121.280 ;
        RECT 257.495 120.780 259.465 121.310 ;
        RECT 278.490 120.780 280.460 121.310 ;
        RECT 283.325 121.330 283.495 121.500 ;
        RECT 283.685 121.330 283.855 121.500 ;
        RECT 284.045 121.330 284.215 121.500 ;
        RECT 284.405 121.330 284.575 121.500 ;
        RECT 284.765 121.330 284.935 121.500 ;
        RECT 285.125 121.330 285.295 121.500 ;
        RECT 330.320 121.330 330.490 121.500 ;
        RECT 330.680 121.330 330.850 121.500 ;
        RECT 331.040 121.330 331.210 121.500 ;
        RECT 331.400 121.330 331.570 121.500 ;
        RECT 331.760 121.330 331.930 121.500 ;
        RECT 332.120 121.330 332.290 121.500 ;
        RECT 205.435 120.280 205.605 120.450 ;
        RECT 205.795 120.280 205.965 120.450 ;
        RECT 206.155 120.280 206.325 120.450 ;
        RECT 206.515 120.280 206.685 120.450 ;
        RECT 206.875 120.280 207.045 120.450 ;
        RECT 207.235 120.280 207.405 120.450 ;
        RECT 252.430 120.280 252.600 120.450 ;
        RECT 252.790 120.280 252.960 120.450 ;
        RECT 253.150 120.280 253.320 120.450 ;
        RECT 253.510 120.280 253.680 120.450 ;
        RECT 253.870 120.280 254.040 120.450 ;
        RECT 254.230 120.280 254.400 120.450 ;
        RECT 283.325 120.500 283.495 120.670 ;
        RECT 283.685 120.500 283.855 120.670 ;
        RECT 284.045 120.500 284.215 120.670 ;
        RECT 284.405 120.500 284.575 120.670 ;
        RECT 284.765 120.500 284.935 120.670 ;
        RECT 285.125 120.500 285.295 120.670 ;
        RECT 330.320 120.500 330.490 120.670 ;
        RECT 330.680 120.500 330.850 120.670 ;
        RECT 331.040 120.500 331.210 120.670 ;
        RECT 331.400 120.500 331.570 120.670 ;
        RECT 331.760 120.500 331.930 120.670 ;
        RECT 332.120 120.500 332.290 120.670 ;
        RECT 205.435 119.450 205.605 119.620 ;
        RECT 205.795 119.450 205.965 119.620 ;
        RECT 206.155 119.450 206.325 119.620 ;
        RECT 206.515 119.450 206.685 119.620 ;
        RECT 206.875 119.450 207.045 119.620 ;
        RECT 207.235 119.450 207.405 119.620 ;
        RECT 252.430 119.450 252.600 119.620 ;
        RECT 252.790 119.450 252.960 119.620 ;
        RECT 253.150 119.450 253.320 119.620 ;
        RECT 253.510 119.450 253.680 119.620 ;
        RECT 253.870 119.450 254.040 119.620 ;
        RECT 254.230 119.450 254.400 119.620 ;
        RECT 257.495 119.610 259.465 120.140 ;
        RECT 278.490 119.610 280.460 120.140 ;
        RECT 283.325 119.670 283.495 119.840 ;
        RECT 283.685 119.670 283.855 119.840 ;
        RECT 284.045 119.670 284.215 119.840 ;
        RECT 284.405 119.670 284.575 119.840 ;
        RECT 284.765 119.670 284.935 119.840 ;
        RECT 285.125 119.670 285.295 119.840 ;
        RECT 330.320 119.670 330.490 119.840 ;
        RECT 330.680 119.670 330.850 119.840 ;
        RECT 331.040 119.670 331.210 119.840 ;
        RECT 331.400 119.670 331.570 119.840 ;
        RECT 331.760 119.670 331.930 119.840 ;
        RECT 332.120 119.670 332.290 119.840 ;
        RECT 205.435 118.620 205.605 118.790 ;
        RECT 205.795 118.620 205.965 118.790 ;
        RECT 206.155 118.620 206.325 118.790 ;
        RECT 206.515 118.620 206.685 118.790 ;
        RECT 206.875 118.620 207.045 118.790 ;
        RECT 207.235 118.620 207.405 118.790 ;
        RECT 252.430 118.620 252.600 118.790 ;
        RECT 252.790 118.620 252.960 118.790 ;
        RECT 253.150 118.620 253.320 118.790 ;
        RECT 253.510 118.620 253.680 118.790 ;
        RECT 253.870 118.620 254.040 118.790 ;
        RECT 254.230 118.620 254.400 118.790 ;
        RECT 257.495 118.440 259.465 118.970 ;
        RECT 278.490 118.440 280.460 118.970 ;
        RECT 283.325 118.840 283.495 119.010 ;
        RECT 283.685 118.840 283.855 119.010 ;
        RECT 284.045 118.840 284.215 119.010 ;
        RECT 284.405 118.840 284.575 119.010 ;
        RECT 284.765 118.840 284.935 119.010 ;
        RECT 285.125 118.840 285.295 119.010 ;
        RECT 330.320 118.840 330.490 119.010 ;
        RECT 330.680 118.840 330.850 119.010 ;
        RECT 331.040 118.840 331.210 119.010 ;
        RECT 331.400 118.840 331.570 119.010 ;
        RECT 331.760 118.840 331.930 119.010 ;
        RECT 332.120 118.840 332.290 119.010 ;
        RECT 205.435 117.790 205.605 117.960 ;
        RECT 205.795 117.790 205.965 117.960 ;
        RECT 206.155 117.790 206.325 117.960 ;
        RECT 206.515 117.790 206.685 117.960 ;
        RECT 206.875 117.790 207.045 117.960 ;
        RECT 207.235 117.790 207.405 117.960 ;
        RECT 252.430 117.790 252.600 117.960 ;
        RECT 252.790 117.790 252.960 117.960 ;
        RECT 253.150 117.790 253.320 117.960 ;
        RECT 253.510 117.790 253.680 117.960 ;
        RECT 253.870 117.790 254.040 117.960 ;
        RECT 254.230 117.790 254.400 117.960 ;
        RECT 283.325 118.010 283.495 118.180 ;
        RECT 283.685 118.010 283.855 118.180 ;
        RECT 284.045 118.010 284.215 118.180 ;
        RECT 284.405 118.010 284.575 118.180 ;
        RECT 284.765 118.010 284.935 118.180 ;
        RECT 285.125 118.010 285.295 118.180 ;
        RECT 330.320 118.010 330.490 118.180 ;
        RECT 330.680 118.010 330.850 118.180 ;
        RECT 331.040 118.010 331.210 118.180 ;
        RECT 331.400 118.010 331.570 118.180 ;
        RECT 331.760 118.010 331.930 118.180 ;
        RECT 332.120 118.010 332.290 118.180 ;
        RECT 257.495 117.270 259.465 117.800 ;
        RECT 205.435 116.960 205.605 117.130 ;
        RECT 205.795 116.960 205.965 117.130 ;
        RECT 206.155 116.960 206.325 117.130 ;
        RECT 206.515 116.960 206.685 117.130 ;
        RECT 206.875 116.960 207.045 117.130 ;
        RECT 207.235 116.960 207.405 117.130 ;
        RECT 278.490 117.270 280.460 117.800 ;
        RECT 252.430 116.960 252.600 117.130 ;
        RECT 252.790 116.960 252.960 117.130 ;
        RECT 253.150 116.960 253.320 117.130 ;
        RECT 253.510 116.960 253.680 117.130 ;
        RECT 253.870 116.960 254.040 117.130 ;
        RECT 254.230 116.960 254.400 117.130 ;
        RECT 283.325 117.180 283.495 117.350 ;
        RECT 283.685 117.180 283.855 117.350 ;
        RECT 284.045 117.180 284.215 117.350 ;
        RECT 284.405 117.180 284.575 117.350 ;
        RECT 284.765 117.180 284.935 117.350 ;
        RECT 285.125 117.180 285.295 117.350 ;
        RECT 330.320 117.180 330.490 117.350 ;
        RECT 330.680 117.180 330.850 117.350 ;
        RECT 331.040 117.180 331.210 117.350 ;
        RECT 331.400 117.180 331.570 117.350 ;
        RECT 331.760 117.180 331.930 117.350 ;
        RECT 332.120 117.180 332.290 117.350 ;
        RECT 205.435 116.130 205.605 116.300 ;
        RECT 205.795 116.130 205.965 116.300 ;
        RECT 206.155 116.130 206.325 116.300 ;
        RECT 206.515 116.130 206.685 116.300 ;
        RECT 206.875 116.130 207.045 116.300 ;
        RECT 207.235 116.130 207.405 116.300 ;
        RECT 252.430 116.130 252.600 116.300 ;
        RECT 252.790 116.130 252.960 116.300 ;
        RECT 253.150 116.130 253.320 116.300 ;
        RECT 253.510 116.130 253.680 116.300 ;
        RECT 253.870 116.130 254.040 116.300 ;
        RECT 254.230 116.130 254.400 116.300 ;
        RECT 257.495 116.100 259.465 116.630 ;
        RECT 278.490 116.100 280.460 116.630 ;
        RECT 283.325 116.350 283.495 116.520 ;
        RECT 283.685 116.350 283.855 116.520 ;
        RECT 284.045 116.350 284.215 116.520 ;
        RECT 284.405 116.350 284.575 116.520 ;
        RECT 284.765 116.350 284.935 116.520 ;
        RECT 285.125 116.350 285.295 116.520 ;
        RECT 330.320 116.350 330.490 116.520 ;
        RECT 330.680 116.350 330.850 116.520 ;
        RECT 331.040 116.350 331.210 116.520 ;
        RECT 331.400 116.350 331.570 116.520 ;
        RECT 331.760 116.350 331.930 116.520 ;
        RECT 332.120 116.350 332.290 116.520 ;
        RECT 205.435 115.300 205.605 115.470 ;
        RECT 205.795 115.300 205.965 115.470 ;
        RECT 206.155 115.300 206.325 115.470 ;
        RECT 206.515 115.300 206.685 115.470 ;
        RECT 206.875 115.300 207.045 115.470 ;
        RECT 207.235 115.300 207.405 115.470 ;
        RECT 252.430 115.300 252.600 115.470 ;
        RECT 252.790 115.300 252.960 115.470 ;
        RECT 253.150 115.300 253.320 115.470 ;
        RECT 253.510 115.300 253.680 115.470 ;
        RECT 253.870 115.300 254.040 115.470 ;
        RECT 254.230 115.300 254.400 115.470 ;
        RECT 257.495 114.930 259.465 115.460 ;
        RECT 278.490 114.930 280.460 115.460 ;
        RECT 283.325 115.520 283.495 115.690 ;
        RECT 283.685 115.520 283.855 115.690 ;
        RECT 284.045 115.520 284.215 115.690 ;
        RECT 284.405 115.520 284.575 115.690 ;
        RECT 284.765 115.520 284.935 115.690 ;
        RECT 285.125 115.520 285.295 115.690 ;
        RECT 330.320 115.520 330.490 115.690 ;
        RECT 330.680 115.520 330.850 115.690 ;
        RECT 331.040 115.520 331.210 115.690 ;
        RECT 331.400 115.520 331.570 115.690 ;
        RECT 331.760 115.520 331.930 115.690 ;
        RECT 332.120 115.520 332.290 115.690 ;
        RECT 205.435 114.470 205.605 114.640 ;
        RECT 205.795 114.470 205.965 114.640 ;
        RECT 206.155 114.470 206.325 114.640 ;
        RECT 206.515 114.470 206.685 114.640 ;
        RECT 206.875 114.470 207.045 114.640 ;
        RECT 207.235 114.470 207.405 114.640 ;
        RECT 252.430 114.470 252.600 114.640 ;
        RECT 252.790 114.470 252.960 114.640 ;
        RECT 253.150 114.470 253.320 114.640 ;
        RECT 253.510 114.470 253.680 114.640 ;
        RECT 253.870 114.470 254.040 114.640 ;
        RECT 254.230 114.470 254.400 114.640 ;
        RECT 283.325 114.690 283.495 114.860 ;
        RECT 283.685 114.690 283.855 114.860 ;
        RECT 284.045 114.690 284.215 114.860 ;
        RECT 284.405 114.690 284.575 114.860 ;
        RECT 284.765 114.690 284.935 114.860 ;
        RECT 285.125 114.690 285.295 114.860 ;
        RECT 330.320 114.690 330.490 114.860 ;
        RECT 330.680 114.690 330.850 114.860 ;
        RECT 331.040 114.690 331.210 114.860 ;
        RECT 331.400 114.690 331.570 114.860 ;
        RECT 331.760 114.690 331.930 114.860 ;
        RECT 332.120 114.690 332.290 114.860 ;
        RECT 205.435 113.640 205.605 113.810 ;
        RECT 205.795 113.640 205.965 113.810 ;
        RECT 206.155 113.640 206.325 113.810 ;
        RECT 206.515 113.640 206.685 113.810 ;
        RECT 206.875 113.640 207.045 113.810 ;
        RECT 207.235 113.640 207.405 113.810 ;
        RECT 252.430 113.640 252.600 113.810 ;
        RECT 252.790 113.640 252.960 113.810 ;
        RECT 253.150 113.640 253.320 113.810 ;
        RECT 253.510 113.640 253.680 113.810 ;
        RECT 253.870 113.640 254.040 113.810 ;
        RECT 254.230 113.640 254.400 113.810 ;
        RECT 257.495 113.760 259.465 114.290 ;
        RECT 278.490 113.760 280.460 114.290 ;
        RECT 283.325 113.860 283.495 114.030 ;
        RECT 283.685 113.860 283.855 114.030 ;
        RECT 284.045 113.860 284.215 114.030 ;
        RECT 284.405 113.860 284.575 114.030 ;
        RECT 284.765 113.860 284.935 114.030 ;
        RECT 285.125 113.860 285.295 114.030 ;
        RECT 330.320 113.860 330.490 114.030 ;
        RECT 330.680 113.860 330.850 114.030 ;
        RECT 331.040 113.860 331.210 114.030 ;
        RECT 331.400 113.860 331.570 114.030 ;
        RECT 331.760 113.860 331.930 114.030 ;
        RECT 332.120 113.860 332.290 114.030 ;
        RECT 205.435 112.810 205.605 112.980 ;
        RECT 205.795 112.810 205.965 112.980 ;
        RECT 206.155 112.810 206.325 112.980 ;
        RECT 206.515 112.810 206.685 112.980 ;
        RECT 206.875 112.810 207.045 112.980 ;
        RECT 207.235 112.810 207.405 112.980 ;
        RECT 252.430 112.810 252.600 112.980 ;
        RECT 252.790 112.810 252.960 112.980 ;
        RECT 253.150 112.810 253.320 112.980 ;
        RECT 253.510 112.810 253.680 112.980 ;
        RECT 253.870 112.810 254.040 112.980 ;
        RECT 254.230 112.810 254.400 112.980 ;
        RECT 257.495 112.590 259.465 113.120 ;
        RECT 278.490 112.590 280.460 113.120 ;
        RECT 283.325 113.030 283.495 113.200 ;
        RECT 283.685 113.030 283.855 113.200 ;
        RECT 284.045 113.030 284.215 113.200 ;
        RECT 284.405 113.030 284.575 113.200 ;
        RECT 284.765 113.030 284.935 113.200 ;
        RECT 285.125 113.030 285.295 113.200 ;
        RECT 330.320 113.030 330.490 113.200 ;
        RECT 330.680 113.030 330.850 113.200 ;
        RECT 331.040 113.030 331.210 113.200 ;
        RECT 331.400 113.030 331.570 113.200 ;
        RECT 331.760 113.030 331.930 113.200 ;
        RECT 332.120 113.030 332.290 113.200 ;
        RECT 205.435 111.980 205.605 112.150 ;
        RECT 205.795 111.980 205.965 112.150 ;
        RECT 206.155 111.980 206.325 112.150 ;
        RECT 206.515 111.980 206.685 112.150 ;
        RECT 206.875 111.980 207.045 112.150 ;
        RECT 207.235 111.980 207.405 112.150 ;
        RECT 252.430 111.980 252.600 112.150 ;
        RECT 252.790 111.980 252.960 112.150 ;
        RECT 253.150 111.980 253.320 112.150 ;
        RECT 253.510 111.980 253.680 112.150 ;
        RECT 253.870 111.980 254.040 112.150 ;
        RECT 254.230 111.980 254.400 112.150 ;
        RECT 283.325 112.200 283.495 112.370 ;
        RECT 283.685 112.200 283.855 112.370 ;
        RECT 284.045 112.200 284.215 112.370 ;
        RECT 284.405 112.200 284.575 112.370 ;
        RECT 284.765 112.200 284.935 112.370 ;
        RECT 285.125 112.200 285.295 112.370 ;
        RECT 330.320 112.200 330.490 112.370 ;
        RECT 330.680 112.200 330.850 112.370 ;
        RECT 331.040 112.200 331.210 112.370 ;
        RECT 331.400 112.200 331.570 112.370 ;
        RECT 331.760 112.200 331.930 112.370 ;
        RECT 332.120 112.200 332.290 112.370 ;
        RECT 257.495 111.420 259.465 111.950 ;
        RECT 205.435 111.150 205.605 111.320 ;
        RECT 205.795 111.150 205.965 111.320 ;
        RECT 206.155 111.150 206.325 111.320 ;
        RECT 206.515 111.150 206.685 111.320 ;
        RECT 206.875 111.150 207.045 111.320 ;
        RECT 207.235 111.150 207.405 111.320 ;
        RECT 278.490 111.420 280.460 111.950 ;
        RECT 283.325 111.370 283.495 111.540 ;
        RECT 283.685 111.370 283.855 111.540 ;
        RECT 284.045 111.370 284.215 111.540 ;
        RECT 284.405 111.370 284.575 111.540 ;
        RECT 284.765 111.370 284.935 111.540 ;
        RECT 285.125 111.370 285.295 111.540 ;
        RECT 252.430 111.150 252.600 111.320 ;
        RECT 252.790 111.150 252.960 111.320 ;
        RECT 253.150 111.150 253.320 111.320 ;
        RECT 253.510 111.150 253.680 111.320 ;
        RECT 253.870 111.150 254.040 111.320 ;
        RECT 254.230 111.150 254.400 111.320 ;
        RECT 330.320 111.370 330.490 111.540 ;
        RECT 330.680 111.370 330.850 111.540 ;
        RECT 331.040 111.370 331.210 111.540 ;
        RECT 331.400 111.370 331.570 111.540 ;
        RECT 331.760 111.370 331.930 111.540 ;
        RECT 332.120 111.370 332.290 111.540 ;
        RECT 205.435 110.320 205.605 110.490 ;
        RECT 205.795 110.320 205.965 110.490 ;
        RECT 206.155 110.320 206.325 110.490 ;
        RECT 206.515 110.320 206.685 110.490 ;
        RECT 206.875 110.320 207.045 110.490 ;
        RECT 207.235 110.320 207.405 110.490 ;
        RECT 252.430 110.320 252.600 110.490 ;
        RECT 252.790 110.320 252.960 110.490 ;
        RECT 253.150 110.320 253.320 110.490 ;
        RECT 253.510 110.320 253.680 110.490 ;
        RECT 253.870 110.320 254.040 110.490 ;
        RECT 254.230 110.320 254.400 110.490 ;
        RECT 257.495 110.250 259.465 110.780 ;
        RECT 278.490 110.250 280.460 110.780 ;
        RECT 283.325 110.540 283.495 110.710 ;
        RECT 283.685 110.540 283.855 110.710 ;
        RECT 284.045 110.540 284.215 110.710 ;
        RECT 284.405 110.540 284.575 110.710 ;
        RECT 284.765 110.540 284.935 110.710 ;
        RECT 285.125 110.540 285.295 110.710 ;
        RECT 330.320 110.540 330.490 110.710 ;
        RECT 330.680 110.540 330.850 110.710 ;
        RECT 331.040 110.540 331.210 110.710 ;
        RECT 331.400 110.540 331.570 110.710 ;
        RECT 331.760 110.540 331.930 110.710 ;
        RECT 332.120 110.540 332.290 110.710 ;
        RECT 205.435 109.490 205.605 109.660 ;
        RECT 205.795 109.490 205.965 109.660 ;
        RECT 206.155 109.490 206.325 109.660 ;
        RECT 206.515 109.490 206.685 109.660 ;
        RECT 206.875 109.490 207.045 109.660 ;
        RECT 207.235 109.490 207.405 109.660 ;
        RECT 283.325 109.710 283.495 109.880 ;
        RECT 283.685 109.710 283.855 109.880 ;
        RECT 284.045 109.710 284.215 109.880 ;
        RECT 284.405 109.710 284.575 109.880 ;
        RECT 284.765 109.710 284.935 109.880 ;
        RECT 285.125 109.710 285.295 109.880 ;
        RECT 252.430 109.490 252.600 109.660 ;
        RECT 252.790 109.490 252.960 109.660 ;
        RECT 253.150 109.490 253.320 109.660 ;
        RECT 253.510 109.490 253.680 109.660 ;
        RECT 253.870 109.490 254.040 109.660 ;
        RECT 254.230 109.490 254.400 109.660 ;
        RECT 257.495 109.080 259.465 109.610 ;
        RECT 330.320 109.710 330.490 109.880 ;
        RECT 330.680 109.710 330.850 109.880 ;
        RECT 331.040 109.710 331.210 109.880 ;
        RECT 331.400 109.710 331.570 109.880 ;
        RECT 331.760 109.710 331.930 109.880 ;
        RECT 332.120 109.710 332.290 109.880 ;
        RECT 278.490 109.080 280.460 109.610 ;
        RECT 205.435 108.660 205.605 108.830 ;
        RECT 205.795 108.660 205.965 108.830 ;
        RECT 206.155 108.660 206.325 108.830 ;
        RECT 206.515 108.660 206.685 108.830 ;
        RECT 206.875 108.660 207.045 108.830 ;
        RECT 207.235 108.660 207.405 108.830 ;
        RECT 252.430 108.660 252.600 108.830 ;
        RECT 252.790 108.660 252.960 108.830 ;
        RECT 253.150 108.660 253.320 108.830 ;
        RECT 253.510 108.660 253.680 108.830 ;
        RECT 253.870 108.660 254.040 108.830 ;
        RECT 254.230 108.660 254.400 108.830 ;
        RECT 283.325 108.880 283.495 109.050 ;
        RECT 283.685 108.880 283.855 109.050 ;
        RECT 284.045 108.880 284.215 109.050 ;
        RECT 284.405 108.880 284.575 109.050 ;
        RECT 284.765 108.880 284.935 109.050 ;
        RECT 285.125 108.880 285.295 109.050 ;
        RECT 330.320 108.880 330.490 109.050 ;
        RECT 330.680 108.880 330.850 109.050 ;
        RECT 331.040 108.880 331.210 109.050 ;
        RECT 331.400 108.880 331.570 109.050 ;
        RECT 331.760 108.880 331.930 109.050 ;
        RECT 332.120 108.880 332.290 109.050 ;
        RECT 205.435 107.830 205.605 108.000 ;
        RECT 205.795 107.830 205.965 108.000 ;
        RECT 206.155 107.830 206.325 108.000 ;
        RECT 206.515 107.830 206.685 108.000 ;
        RECT 206.875 107.830 207.045 108.000 ;
        RECT 207.235 107.830 207.405 108.000 ;
        RECT 252.430 107.830 252.600 108.000 ;
        RECT 252.790 107.830 252.960 108.000 ;
        RECT 253.150 107.830 253.320 108.000 ;
        RECT 253.510 107.830 253.680 108.000 ;
        RECT 253.870 107.830 254.040 108.000 ;
        RECT 254.230 107.830 254.400 108.000 ;
        RECT 257.495 107.910 259.465 108.440 ;
        RECT 278.490 107.910 280.460 108.440 ;
        RECT 283.325 108.050 283.495 108.220 ;
        RECT 283.685 108.050 283.855 108.220 ;
        RECT 284.045 108.050 284.215 108.220 ;
        RECT 284.405 108.050 284.575 108.220 ;
        RECT 284.765 108.050 284.935 108.220 ;
        RECT 285.125 108.050 285.295 108.220 ;
        RECT 330.320 108.050 330.490 108.220 ;
        RECT 330.680 108.050 330.850 108.220 ;
        RECT 331.040 108.050 331.210 108.220 ;
        RECT 331.400 108.050 331.570 108.220 ;
        RECT 331.760 108.050 331.930 108.220 ;
        RECT 332.120 108.050 332.290 108.220 ;
        RECT 205.435 107.000 205.605 107.170 ;
        RECT 205.795 107.000 205.965 107.170 ;
        RECT 206.155 107.000 206.325 107.170 ;
        RECT 206.515 107.000 206.685 107.170 ;
        RECT 206.875 107.000 207.045 107.170 ;
        RECT 207.235 107.000 207.405 107.170 ;
        RECT 252.430 107.000 252.600 107.170 ;
        RECT 252.790 107.000 252.960 107.170 ;
        RECT 253.150 107.000 253.320 107.170 ;
        RECT 253.510 107.000 253.680 107.170 ;
        RECT 253.870 107.000 254.040 107.170 ;
        RECT 254.230 107.000 254.400 107.170 ;
        RECT 257.495 106.740 259.465 107.270 ;
        RECT 278.490 106.740 280.460 107.270 ;
        RECT 283.325 107.220 283.495 107.390 ;
        RECT 283.685 107.220 283.855 107.390 ;
        RECT 284.045 107.220 284.215 107.390 ;
        RECT 284.405 107.220 284.575 107.390 ;
        RECT 284.765 107.220 284.935 107.390 ;
        RECT 285.125 107.220 285.295 107.390 ;
        RECT 330.320 107.220 330.490 107.390 ;
        RECT 330.680 107.220 330.850 107.390 ;
        RECT 331.040 107.220 331.210 107.390 ;
        RECT 331.400 107.220 331.570 107.390 ;
        RECT 331.760 107.220 331.930 107.390 ;
        RECT 332.120 107.220 332.290 107.390 ;
        RECT 205.435 106.170 205.605 106.340 ;
        RECT 205.795 106.170 205.965 106.340 ;
        RECT 206.155 106.170 206.325 106.340 ;
        RECT 206.515 106.170 206.685 106.340 ;
        RECT 206.875 106.170 207.045 106.340 ;
        RECT 207.235 106.170 207.405 106.340 ;
        RECT 252.430 106.170 252.600 106.340 ;
        RECT 252.790 106.170 252.960 106.340 ;
        RECT 253.150 106.170 253.320 106.340 ;
        RECT 253.510 106.170 253.680 106.340 ;
        RECT 253.870 106.170 254.040 106.340 ;
        RECT 254.230 106.170 254.400 106.340 ;
        RECT 283.325 106.390 283.495 106.560 ;
        RECT 283.685 106.390 283.855 106.560 ;
        RECT 284.045 106.390 284.215 106.560 ;
        RECT 284.405 106.390 284.575 106.560 ;
        RECT 284.765 106.390 284.935 106.560 ;
        RECT 285.125 106.390 285.295 106.560 ;
        RECT 330.320 106.390 330.490 106.560 ;
        RECT 330.680 106.390 330.850 106.560 ;
        RECT 331.040 106.390 331.210 106.560 ;
        RECT 331.400 106.390 331.570 106.560 ;
        RECT 331.760 106.390 331.930 106.560 ;
        RECT 332.120 106.390 332.290 106.560 ;
        RECT 205.435 105.340 205.605 105.510 ;
        RECT 205.795 105.340 205.965 105.510 ;
        RECT 206.155 105.340 206.325 105.510 ;
        RECT 206.515 105.340 206.685 105.510 ;
        RECT 206.875 105.340 207.045 105.510 ;
        RECT 207.235 105.340 207.405 105.510 ;
        RECT 252.430 105.340 252.600 105.510 ;
        RECT 252.790 105.340 252.960 105.510 ;
        RECT 253.150 105.340 253.320 105.510 ;
        RECT 253.510 105.340 253.680 105.510 ;
        RECT 253.870 105.340 254.040 105.510 ;
        RECT 254.230 105.340 254.400 105.510 ;
        RECT 257.495 105.570 259.465 106.100 ;
        RECT 278.490 105.570 280.460 106.100 ;
        RECT 283.325 105.560 283.495 105.730 ;
        RECT 283.685 105.560 283.855 105.730 ;
        RECT 284.045 105.560 284.215 105.730 ;
        RECT 284.405 105.560 284.575 105.730 ;
        RECT 284.765 105.560 284.935 105.730 ;
        RECT 285.125 105.560 285.295 105.730 ;
        RECT 330.320 105.560 330.490 105.730 ;
        RECT 330.680 105.560 330.850 105.730 ;
        RECT 331.040 105.560 331.210 105.730 ;
        RECT 331.400 105.560 331.570 105.730 ;
        RECT 331.760 105.560 331.930 105.730 ;
        RECT 332.120 105.560 332.290 105.730 ;
        RECT 205.435 104.510 205.605 104.680 ;
        RECT 205.795 104.510 205.965 104.680 ;
        RECT 206.155 104.510 206.325 104.680 ;
        RECT 206.515 104.510 206.685 104.680 ;
        RECT 206.875 104.510 207.045 104.680 ;
        RECT 207.235 104.510 207.405 104.680 ;
        RECT 252.430 104.510 252.600 104.680 ;
        RECT 252.790 104.510 252.960 104.680 ;
        RECT 253.150 104.510 253.320 104.680 ;
        RECT 253.510 104.510 253.680 104.680 ;
        RECT 253.870 104.510 254.040 104.680 ;
        RECT 254.230 104.510 254.400 104.680 ;
        RECT 257.495 104.400 259.465 104.930 ;
        RECT 278.490 104.400 280.460 104.930 ;
        RECT 283.325 104.730 283.495 104.900 ;
        RECT 283.685 104.730 283.855 104.900 ;
        RECT 284.045 104.730 284.215 104.900 ;
        RECT 284.405 104.730 284.575 104.900 ;
        RECT 284.765 104.730 284.935 104.900 ;
        RECT 285.125 104.730 285.295 104.900 ;
        RECT 330.320 104.730 330.490 104.900 ;
        RECT 330.680 104.730 330.850 104.900 ;
        RECT 331.040 104.730 331.210 104.900 ;
        RECT 331.400 104.730 331.570 104.900 ;
        RECT 331.760 104.730 331.930 104.900 ;
        RECT 332.120 104.730 332.290 104.900 ;
        RECT 205.435 103.680 205.605 103.850 ;
        RECT 205.795 103.680 205.965 103.850 ;
        RECT 206.155 103.680 206.325 103.850 ;
        RECT 206.515 103.680 206.685 103.850 ;
        RECT 206.875 103.680 207.045 103.850 ;
        RECT 207.235 103.680 207.405 103.850 ;
        RECT 252.430 103.680 252.600 103.850 ;
        RECT 252.790 103.680 252.960 103.850 ;
        RECT 253.150 103.680 253.320 103.850 ;
        RECT 253.510 103.680 253.680 103.850 ;
        RECT 253.870 103.680 254.040 103.850 ;
        RECT 254.230 103.680 254.400 103.850 ;
        RECT 283.325 103.900 283.495 104.070 ;
        RECT 283.685 103.900 283.855 104.070 ;
        RECT 284.045 103.900 284.215 104.070 ;
        RECT 284.405 103.900 284.575 104.070 ;
        RECT 284.765 103.900 284.935 104.070 ;
        RECT 285.125 103.900 285.295 104.070 ;
        RECT 257.495 103.230 259.465 103.760 ;
        RECT 330.320 103.900 330.490 104.070 ;
        RECT 330.680 103.900 330.850 104.070 ;
        RECT 331.040 103.900 331.210 104.070 ;
        RECT 331.400 103.900 331.570 104.070 ;
        RECT 331.760 103.900 331.930 104.070 ;
        RECT 332.120 103.900 332.290 104.070 ;
        RECT 278.490 103.230 280.460 103.760 ;
        RECT 205.435 102.850 205.605 103.020 ;
        RECT 205.795 102.850 205.965 103.020 ;
        RECT 206.155 102.850 206.325 103.020 ;
        RECT 206.515 102.850 206.685 103.020 ;
        RECT 206.875 102.850 207.045 103.020 ;
        RECT 207.235 102.850 207.405 103.020 ;
        RECT 252.430 102.850 252.600 103.020 ;
        RECT 252.790 102.850 252.960 103.020 ;
        RECT 253.150 102.850 253.320 103.020 ;
        RECT 253.510 102.850 253.680 103.020 ;
        RECT 253.870 102.850 254.040 103.020 ;
        RECT 254.230 102.850 254.400 103.020 ;
        RECT 283.325 103.070 283.495 103.240 ;
        RECT 283.685 103.070 283.855 103.240 ;
        RECT 284.045 103.070 284.215 103.240 ;
        RECT 284.405 103.070 284.575 103.240 ;
        RECT 284.765 103.070 284.935 103.240 ;
        RECT 285.125 103.070 285.295 103.240 ;
        RECT 330.320 103.070 330.490 103.240 ;
        RECT 330.680 103.070 330.850 103.240 ;
        RECT 331.040 103.070 331.210 103.240 ;
        RECT 331.400 103.070 331.570 103.240 ;
        RECT 331.760 103.070 331.930 103.240 ;
        RECT 332.120 103.070 332.290 103.240 ;
        RECT 205.435 102.020 205.605 102.190 ;
        RECT 205.795 102.020 205.965 102.190 ;
        RECT 206.155 102.020 206.325 102.190 ;
        RECT 206.515 102.020 206.685 102.190 ;
        RECT 206.875 102.020 207.045 102.190 ;
        RECT 207.235 102.020 207.405 102.190 ;
        RECT 252.430 102.020 252.600 102.190 ;
        RECT 252.790 102.020 252.960 102.190 ;
        RECT 253.150 102.020 253.320 102.190 ;
        RECT 253.510 102.020 253.680 102.190 ;
        RECT 253.870 102.020 254.040 102.190 ;
        RECT 254.230 102.020 254.400 102.190 ;
        RECT 283.325 102.240 283.495 102.410 ;
        RECT 283.685 102.240 283.855 102.410 ;
        RECT 284.045 102.240 284.215 102.410 ;
        RECT 284.405 102.240 284.575 102.410 ;
        RECT 284.765 102.240 284.935 102.410 ;
        RECT 285.125 102.240 285.295 102.410 ;
        RECT 330.320 102.240 330.490 102.410 ;
        RECT 330.680 102.240 330.850 102.410 ;
        RECT 331.040 102.240 331.210 102.410 ;
        RECT 331.400 102.240 331.570 102.410 ;
        RECT 331.760 102.240 331.930 102.410 ;
        RECT 332.120 102.240 332.290 102.410 ;
        RECT 205.435 101.190 205.605 101.360 ;
        RECT 205.795 101.190 205.965 101.360 ;
        RECT 206.155 101.190 206.325 101.360 ;
        RECT 206.515 101.190 206.685 101.360 ;
        RECT 206.875 101.190 207.045 101.360 ;
        RECT 207.235 101.190 207.405 101.360 ;
        RECT 252.430 101.190 252.600 101.360 ;
        RECT 252.790 101.190 252.960 101.360 ;
        RECT 253.150 101.190 253.320 101.360 ;
        RECT 253.510 101.190 253.680 101.360 ;
        RECT 253.870 101.190 254.040 101.360 ;
        RECT 254.230 101.190 254.400 101.360 ;
        RECT 283.325 101.410 283.495 101.580 ;
        RECT 283.685 101.410 283.855 101.580 ;
        RECT 284.045 101.410 284.215 101.580 ;
        RECT 284.405 101.410 284.575 101.580 ;
        RECT 284.765 101.410 284.935 101.580 ;
        RECT 285.125 101.410 285.295 101.580 ;
        RECT 330.320 101.410 330.490 101.580 ;
        RECT 330.680 101.410 330.850 101.580 ;
        RECT 331.040 101.410 331.210 101.580 ;
        RECT 331.400 101.410 331.570 101.580 ;
        RECT 331.760 101.410 331.930 101.580 ;
        RECT 332.120 101.410 332.290 101.580 ;
        RECT 205.435 100.360 205.605 100.530 ;
        RECT 205.795 100.360 205.965 100.530 ;
        RECT 206.155 100.360 206.325 100.530 ;
        RECT 206.515 100.360 206.685 100.530 ;
        RECT 206.875 100.360 207.045 100.530 ;
        RECT 207.235 100.360 207.405 100.530 ;
        RECT 252.430 100.360 252.600 100.530 ;
        RECT 252.790 100.360 252.960 100.530 ;
        RECT 253.150 100.360 253.320 100.530 ;
        RECT 253.510 100.360 253.680 100.530 ;
        RECT 253.870 100.360 254.040 100.530 ;
        RECT 254.230 100.360 254.400 100.530 ;
        RECT 283.325 100.580 283.495 100.750 ;
        RECT 283.685 100.580 283.855 100.750 ;
        RECT 284.045 100.580 284.215 100.750 ;
        RECT 284.405 100.580 284.575 100.750 ;
        RECT 284.765 100.580 284.935 100.750 ;
        RECT 285.125 100.580 285.295 100.750 ;
        RECT 330.320 100.580 330.490 100.750 ;
        RECT 330.680 100.580 330.850 100.750 ;
        RECT 331.040 100.580 331.210 100.750 ;
        RECT 331.400 100.580 331.570 100.750 ;
        RECT 331.760 100.580 331.930 100.750 ;
        RECT 332.120 100.580 332.290 100.750 ;
        RECT 205.435 99.530 205.605 99.700 ;
        RECT 205.795 99.530 205.965 99.700 ;
        RECT 206.155 99.530 206.325 99.700 ;
        RECT 206.515 99.530 206.685 99.700 ;
        RECT 206.875 99.530 207.045 99.700 ;
        RECT 207.235 99.530 207.405 99.700 ;
        RECT 252.430 99.530 252.600 99.700 ;
        RECT 252.790 99.530 252.960 99.700 ;
        RECT 253.150 99.530 253.320 99.700 ;
        RECT 253.510 99.530 253.680 99.700 ;
        RECT 253.870 99.530 254.040 99.700 ;
        RECT 254.230 99.530 254.400 99.700 ;
        RECT 283.325 99.750 283.495 99.920 ;
        RECT 283.685 99.750 283.855 99.920 ;
        RECT 284.045 99.750 284.215 99.920 ;
        RECT 284.405 99.750 284.575 99.920 ;
        RECT 284.765 99.750 284.935 99.920 ;
        RECT 285.125 99.750 285.295 99.920 ;
        RECT 330.320 99.750 330.490 99.920 ;
        RECT 330.680 99.750 330.850 99.920 ;
        RECT 331.040 99.750 331.210 99.920 ;
        RECT 331.400 99.750 331.570 99.920 ;
        RECT 331.760 99.750 331.930 99.920 ;
        RECT 332.120 99.750 332.290 99.920 ;
        RECT 270.600 99.180 270.770 99.350 ;
        RECT 273.290 99.180 273.460 99.350 ;
        RECT 205.435 98.700 205.605 98.870 ;
        RECT 205.795 98.700 205.965 98.870 ;
        RECT 206.155 98.700 206.325 98.870 ;
        RECT 206.515 98.700 206.685 98.870 ;
        RECT 206.875 98.700 207.045 98.870 ;
        RECT 207.235 98.700 207.405 98.870 ;
        RECT 252.430 98.700 252.600 98.870 ;
        RECT 252.790 98.700 252.960 98.870 ;
        RECT 253.150 98.700 253.320 98.870 ;
        RECT 253.510 98.700 253.680 98.870 ;
        RECT 253.870 98.700 254.040 98.870 ;
        RECT 254.230 98.700 254.400 98.870 ;
        RECT 266.310 98.700 266.480 98.870 ;
        RECT 270.115 98.785 270.285 98.955 ;
        RECT 273.775 98.785 273.945 98.955 ;
        RECT 283.325 98.920 283.495 99.090 ;
        RECT 283.685 98.920 283.855 99.090 ;
        RECT 284.045 98.920 284.215 99.090 ;
        RECT 284.405 98.920 284.575 99.090 ;
        RECT 284.765 98.920 284.935 99.090 ;
        RECT 285.125 98.920 285.295 99.090 ;
        RECT 330.320 98.920 330.490 99.090 ;
        RECT 330.680 98.920 330.850 99.090 ;
        RECT 331.040 98.920 331.210 99.090 ;
        RECT 331.400 98.920 331.570 99.090 ;
        RECT 331.760 98.920 331.930 99.090 ;
        RECT 332.120 98.920 332.290 99.090 ;
        RECT 266.840 98.305 267.010 98.475 ;
        RECT 270.600 98.390 270.770 98.560 ;
        RECT 205.435 97.870 205.605 98.040 ;
        RECT 205.795 97.870 205.965 98.040 ;
        RECT 206.155 97.870 206.325 98.040 ;
        RECT 206.515 97.870 206.685 98.040 ;
        RECT 206.875 97.870 207.045 98.040 ;
        RECT 207.235 97.870 207.405 98.040 ;
        RECT 252.430 97.870 252.600 98.040 ;
        RECT 252.790 97.870 252.960 98.040 ;
        RECT 253.150 97.870 253.320 98.040 ;
        RECT 253.510 97.870 253.680 98.040 ;
        RECT 253.870 97.870 254.040 98.040 ;
        RECT 254.230 97.870 254.400 98.040 ;
        RECT 283.325 98.090 283.495 98.260 ;
        RECT 283.685 98.090 283.855 98.260 ;
        RECT 284.045 98.090 284.215 98.260 ;
        RECT 284.405 98.090 284.575 98.260 ;
        RECT 284.765 98.090 284.935 98.260 ;
        RECT 285.125 98.090 285.295 98.260 ;
        RECT 330.320 98.090 330.490 98.260 ;
        RECT 330.680 98.090 330.850 98.260 ;
        RECT 331.040 98.090 331.210 98.260 ;
        RECT 331.400 98.090 331.570 98.260 ;
        RECT 331.760 98.090 331.930 98.260 ;
        RECT 332.120 98.090 332.290 98.260 ;
        RECT 205.435 97.040 205.605 97.210 ;
        RECT 205.795 97.040 205.965 97.210 ;
        RECT 206.155 97.040 206.325 97.210 ;
        RECT 206.515 97.040 206.685 97.210 ;
        RECT 206.875 97.040 207.045 97.210 ;
        RECT 207.235 97.040 207.405 97.210 ;
        RECT 252.430 97.040 252.600 97.210 ;
        RECT 252.790 97.040 252.960 97.210 ;
        RECT 253.150 97.040 253.320 97.210 ;
        RECT 253.510 97.040 253.680 97.210 ;
        RECT 253.870 97.040 254.040 97.210 ;
        RECT 254.230 97.040 254.400 97.210 ;
        RECT 283.325 97.260 283.495 97.430 ;
        RECT 283.685 97.260 283.855 97.430 ;
        RECT 284.045 97.260 284.215 97.430 ;
        RECT 284.405 97.260 284.575 97.430 ;
        RECT 284.765 97.260 284.935 97.430 ;
        RECT 285.125 97.260 285.295 97.430 ;
        RECT 330.320 97.260 330.490 97.430 ;
        RECT 330.680 97.260 330.850 97.430 ;
        RECT 331.040 97.260 331.210 97.430 ;
        RECT 331.400 97.260 331.570 97.430 ;
        RECT 331.760 97.260 331.930 97.430 ;
        RECT 332.120 97.260 332.290 97.430 ;
        RECT 205.435 96.210 205.605 96.380 ;
        RECT 205.795 96.210 205.965 96.380 ;
        RECT 206.155 96.210 206.325 96.380 ;
        RECT 206.515 96.210 206.685 96.380 ;
        RECT 206.875 96.210 207.045 96.380 ;
        RECT 207.235 96.210 207.405 96.380 ;
        RECT 270.600 96.400 270.770 96.570 ;
        RECT 273.290 96.400 273.460 96.570 ;
        RECT 283.325 96.430 283.495 96.600 ;
        RECT 283.685 96.430 283.855 96.600 ;
        RECT 284.045 96.430 284.215 96.600 ;
        RECT 284.405 96.430 284.575 96.600 ;
        RECT 284.765 96.430 284.935 96.600 ;
        RECT 285.125 96.430 285.295 96.600 ;
        RECT 252.430 96.210 252.600 96.380 ;
        RECT 252.790 96.210 252.960 96.380 ;
        RECT 253.150 96.210 253.320 96.380 ;
        RECT 253.510 96.210 253.680 96.380 ;
        RECT 253.870 96.210 254.040 96.380 ;
        RECT 254.230 96.210 254.400 96.380 ;
        RECT 330.320 96.430 330.490 96.600 ;
        RECT 330.680 96.430 330.850 96.600 ;
        RECT 331.040 96.430 331.210 96.600 ;
        RECT 331.400 96.430 331.570 96.600 ;
        RECT 331.760 96.430 331.930 96.600 ;
        RECT 332.120 96.430 332.290 96.600 ;
        RECT 270.115 96.005 270.285 96.175 ;
        RECT 273.775 96.005 273.945 96.175 ;
        RECT 205.435 95.380 205.605 95.550 ;
        RECT 205.795 95.380 205.965 95.550 ;
        RECT 206.155 95.380 206.325 95.550 ;
        RECT 206.515 95.380 206.685 95.550 ;
        RECT 206.875 95.380 207.045 95.550 ;
        RECT 207.235 95.380 207.405 95.550 ;
        RECT 266.310 95.620 266.480 95.790 ;
        RECT 270.600 95.610 270.770 95.780 ;
        RECT 283.325 95.600 283.495 95.770 ;
        RECT 283.685 95.600 283.855 95.770 ;
        RECT 284.045 95.600 284.215 95.770 ;
        RECT 284.405 95.600 284.575 95.770 ;
        RECT 284.765 95.600 284.935 95.770 ;
        RECT 285.125 95.600 285.295 95.770 ;
        RECT 252.430 95.380 252.600 95.550 ;
        RECT 252.790 95.380 252.960 95.550 ;
        RECT 253.150 95.380 253.320 95.550 ;
        RECT 253.510 95.380 253.680 95.550 ;
        RECT 253.870 95.380 254.040 95.550 ;
        RECT 254.230 95.380 254.400 95.550 ;
        RECT 262.750 95.225 262.920 95.395 ;
        RECT 330.320 95.600 330.490 95.770 ;
        RECT 330.680 95.600 330.850 95.770 ;
        RECT 331.040 95.600 331.210 95.770 ;
        RECT 331.400 95.600 331.570 95.770 ;
        RECT 331.760 95.600 331.930 95.770 ;
        RECT 332.120 95.600 332.290 95.770 ;
        RECT 266.840 95.225 267.010 95.395 ;
        RECT 263.280 94.830 263.450 95.000 ;
        RECT 266.310 94.830 266.480 95.000 ;
        RECT 205.435 94.550 205.605 94.720 ;
        RECT 205.795 94.550 205.965 94.720 ;
        RECT 206.155 94.550 206.325 94.720 ;
        RECT 206.515 94.550 206.685 94.720 ;
        RECT 206.875 94.550 207.045 94.720 ;
        RECT 207.235 94.550 207.405 94.720 ;
        RECT 252.430 94.550 252.600 94.720 ;
        RECT 252.790 94.550 252.960 94.720 ;
        RECT 253.150 94.550 253.320 94.720 ;
        RECT 253.510 94.550 253.680 94.720 ;
        RECT 253.870 94.550 254.040 94.720 ;
        RECT 254.230 94.550 254.400 94.720 ;
        RECT 283.325 94.770 283.495 94.940 ;
        RECT 283.685 94.770 283.855 94.940 ;
        RECT 284.045 94.770 284.215 94.940 ;
        RECT 284.405 94.770 284.575 94.940 ;
        RECT 284.765 94.770 284.935 94.940 ;
        RECT 285.125 94.770 285.295 94.940 ;
        RECT 330.320 94.770 330.490 94.940 ;
        RECT 330.680 94.770 330.850 94.940 ;
        RECT 331.040 94.770 331.210 94.940 ;
        RECT 331.400 94.770 331.570 94.940 ;
        RECT 331.760 94.770 331.930 94.940 ;
        RECT 332.120 94.770 332.290 94.940 ;
        RECT 205.435 93.720 205.605 93.890 ;
        RECT 205.795 93.720 205.965 93.890 ;
        RECT 206.155 93.720 206.325 93.890 ;
        RECT 206.515 93.720 206.685 93.890 ;
        RECT 206.875 93.720 207.045 93.890 ;
        RECT 207.235 93.720 207.405 93.890 ;
        RECT 252.430 93.720 252.600 93.890 ;
        RECT 252.790 93.720 252.960 93.890 ;
        RECT 253.150 93.720 253.320 93.890 ;
        RECT 253.510 93.720 253.680 93.890 ;
        RECT 253.870 93.720 254.040 93.890 ;
        RECT 254.230 93.720 254.400 93.890 ;
        RECT 283.325 93.940 283.495 94.110 ;
        RECT 283.685 93.940 283.855 94.110 ;
        RECT 284.045 93.940 284.215 94.110 ;
        RECT 284.405 93.940 284.575 94.110 ;
        RECT 284.765 93.940 284.935 94.110 ;
        RECT 285.125 93.940 285.295 94.110 ;
        RECT 330.320 93.940 330.490 94.110 ;
        RECT 330.680 93.940 330.850 94.110 ;
        RECT 331.040 93.940 331.210 94.110 ;
        RECT 331.400 93.940 331.570 94.110 ;
        RECT 331.760 93.940 331.930 94.110 ;
        RECT 332.120 93.940 332.290 94.110 ;
        RECT 270.600 93.620 270.770 93.790 ;
        RECT 273.290 93.620 273.460 93.790 ;
        RECT 276.920 93.610 277.090 93.780 ;
        RECT 270.115 93.225 270.285 93.395 ;
        RECT 205.435 92.890 205.605 93.060 ;
        RECT 205.795 92.890 205.965 93.060 ;
        RECT 206.155 92.890 206.325 93.060 ;
        RECT 206.515 92.890 206.685 93.060 ;
        RECT 206.875 92.890 207.045 93.060 ;
        RECT 207.235 92.890 207.405 93.060 ;
        RECT 273.775 93.225 273.945 93.395 ;
        RECT 277.405 93.215 277.575 93.385 ;
        RECT 252.430 92.890 252.600 93.060 ;
        RECT 252.790 92.890 252.960 93.060 ;
        RECT 253.150 92.890 253.320 93.060 ;
        RECT 253.510 92.890 253.680 93.060 ;
        RECT 253.870 92.890 254.040 93.060 ;
        RECT 254.230 92.890 254.400 93.060 ;
        RECT 283.325 93.110 283.495 93.280 ;
        RECT 283.685 93.110 283.855 93.280 ;
        RECT 284.045 93.110 284.215 93.280 ;
        RECT 284.405 93.110 284.575 93.280 ;
        RECT 284.765 93.110 284.935 93.280 ;
        RECT 285.125 93.110 285.295 93.280 ;
        RECT 330.320 93.110 330.490 93.280 ;
        RECT 330.680 93.110 330.850 93.280 ;
        RECT 331.040 93.110 331.210 93.280 ;
        RECT 331.400 93.110 331.570 93.280 ;
        RECT 331.760 93.110 331.930 93.280 ;
        RECT 332.120 93.110 332.290 93.280 ;
        RECT 270.600 92.830 270.770 93.000 ;
        RECT 266.310 92.540 266.480 92.710 ;
        RECT 205.435 92.060 205.605 92.230 ;
        RECT 205.795 92.060 205.965 92.230 ;
        RECT 206.155 92.060 206.325 92.230 ;
        RECT 206.515 92.060 206.685 92.230 ;
        RECT 206.875 92.060 207.045 92.230 ;
        RECT 207.235 92.060 207.405 92.230 ;
        RECT 252.430 92.060 252.600 92.230 ;
        RECT 252.790 92.060 252.960 92.230 ;
        RECT 253.150 92.060 253.320 92.230 ;
        RECT 253.510 92.060 253.680 92.230 ;
        RECT 253.870 92.060 254.040 92.230 ;
        RECT 254.230 92.060 254.400 92.230 ;
        RECT 262.750 92.145 262.920 92.315 ;
        RECT 266.840 92.145 267.010 92.315 ;
        RECT 283.325 92.280 283.495 92.450 ;
        RECT 283.685 92.280 283.855 92.450 ;
        RECT 284.045 92.280 284.215 92.450 ;
        RECT 284.405 92.280 284.575 92.450 ;
        RECT 284.765 92.280 284.935 92.450 ;
        RECT 285.125 92.280 285.295 92.450 ;
        RECT 330.320 92.280 330.490 92.450 ;
        RECT 330.680 92.280 330.850 92.450 ;
        RECT 331.040 92.280 331.210 92.450 ;
        RECT 331.400 92.280 331.570 92.450 ;
        RECT 331.760 92.280 331.930 92.450 ;
        RECT 332.120 92.280 332.290 92.450 ;
        RECT 263.280 91.750 263.450 91.920 ;
        RECT 266.310 91.750 266.480 91.920 ;
        RECT 205.435 91.230 205.605 91.400 ;
        RECT 205.795 91.230 205.965 91.400 ;
        RECT 206.155 91.230 206.325 91.400 ;
        RECT 206.515 91.230 206.685 91.400 ;
        RECT 206.875 91.230 207.045 91.400 ;
        RECT 207.235 91.230 207.405 91.400 ;
        RECT 252.430 91.230 252.600 91.400 ;
        RECT 252.790 91.230 252.960 91.400 ;
        RECT 253.150 91.230 253.320 91.400 ;
        RECT 253.510 91.230 253.680 91.400 ;
        RECT 253.870 91.230 254.040 91.400 ;
        RECT 254.230 91.230 254.400 91.400 ;
        RECT 283.325 91.450 283.495 91.620 ;
        RECT 283.685 91.450 283.855 91.620 ;
        RECT 284.045 91.450 284.215 91.620 ;
        RECT 284.405 91.450 284.575 91.620 ;
        RECT 284.765 91.450 284.935 91.620 ;
        RECT 285.125 91.450 285.295 91.620 ;
        RECT 330.320 91.450 330.490 91.620 ;
        RECT 330.680 91.450 330.850 91.620 ;
        RECT 331.040 91.450 331.210 91.620 ;
        RECT 331.400 91.450 331.570 91.620 ;
        RECT 331.760 91.450 331.930 91.620 ;
        RECT 332.120 91.450 332.290 91.620 ;
        RECT 270.600 90.840 270.770 91.010 ;
        RECT 273.290 90.840 273.460 91.010 ;
        RECT 205.435 90.400 205.605 90.570 ;
        RECT 205.795 90.400 205.965 90.570 ;
        RECT 206.155 90.400 206.325 90.570 ;
        RECT 206.515 90.400 206.685 90.570 ;
        RECT 206.875 90.400 207.045 90.570 ;
        RECT 207.235 90.400 207.405 90.570 ;
        RECT 252.430 90.400 252.600 90.570 ;
        RECT 252.790 90.400 252.960 90.570 ;
        RECT 253.150 90.400 253.320 90.570 ;
        RECT 253.510 90.400 253.680 90.570 ;
        RECT 253.870 90.400 254.040 90.570 ;
        RECT 254.230 90.400 254.400 90.570 ;
        RECT 273.775 90.445 273.945 90.615 ;
        RECT 277.405 90.435 277.575 90.605 ;
        RECT 283.325 90.620 283.495 90.790 ;
        RECT 283.685 90.620 283.855 90.790 ;
        RECT 284.045 90.620 284.215 90.790 ;
        RECT 284.405 90.620 284.575 90.790 ;
        RECT 284.765 90.620 284.935 90.790 ;
        RECT 285.125 90.620 285.295 90.790 ;
        RECT 330.320 90.620 330.490 90.790 ;
        RECT 330.680 90.620 330.850 90.790 ;
        RECT 331.040 90.620 331.210 90.790 ;
        RECT 331.400 90.620 331.570 90.790 ;
        RECT 331.760 90.620 331.930 90.790 ;
        RECT 332.120 90.620 332.290 90.790 ;
        RECT 270.600 90.050 270.770 90.220 ;
        RECT 205.435 89.570 205.605 89.740 ;
        RECT 205.795 89.570 205.965 89.740 ;
        RECT 206.155 89.570 206.325 89.740 ;
        RECT 206.515 89.570 206.685 89.740 ;
        RECT 206.875 89.570 207.045 89.740 ;
        RECT 207.235 89.570 207.405 89.740 ;
        RECT 252.430 89.570 252.600 89.740 ;
        RECT 252.790 89.570 252.960 89.740 ;
        RECT 253.150 89.570 253.320 89.740 ;
        RECT 253.510 89.570 253.680 89.740 ;
        RECT 253.870 89.570 254.040 89.740 ;
        RECT 254.230 89.570 254.400 89.740 ;
        RECT 283.325 89.790 283.495 89.960 ;
        RECT 283.685 89.790 283.855 89.960 ;
        RECT 284.045 89.790 284.215 89.960 ;
        RECT 284.405 89.790 284.575 89.960 ;
        RECT 284.765 89.790 284.935 89.960 ;
        RECT 285.125 89.790 285.295 89.960 ;
        RECT 330.320 89.790 330.490 89.960 ;
        RECT 330.680 89.790 330.850 89.960 ;
        RECT 331.040 89.790 331.210 89.960 ;
        RECT 331.400 89.790 331.570 89.960 ;
        RECT 331.760 89.790 331.930 89.960 ;
        RECT 332.120 89.790 332.290 89.960 ;
        RECT 266.310 89.460 266.480 89.630 ;
        RECT 262.750 89.065 262.920 89.235 ;
        RECT 205.435 88.740 205.605 88.910 ;
        RECT 205.795 88.740 205.965 88.910 ;
        RECT 206.155 88.740 206.325 88.910 ;
        RECT 206.515 88.740 206.685 88.910 ;
        RECT 206.875 88.740 207.045 88.910 ;
        RECT 207.235 88.740 207.405 88.910 ;
        RECT 252.430 88.740 252.600 88.910 ;
        RECT 252.790 88.740 252.960 88.910 ;
        RECT 253.150 88.740 253.320 88.910 ;
        RECT 253.510 88.740 253.680 88.910 ;
        RECT 253.870 88.740 254.040 88.910 ;
        RECT 254.230 88.740 254.400 88.910 ;
        RECT 283.325 88.960 283.495 89.130 ;
        RECT 283.685 88.960 283.855 89.130 ;
        RECT 284.045 88.960 284.215 89.130 ;
        RECT 284.405 88.960 284.575 89.130 ;
        RECT 284.765 88.960 284.935 89.130 ;
        RECT 285.125 88.960 285.295 89.130 ;
        RECT 330.320 88.960 330.490 89.130 ;
        RECT 330.680 88.960 330.850 89.130 ;
        RECT 331.040 88.960 331.210 89.130 ;
        RECT 331.400 88.960 331.570 89.130 ;
        RECT 331.760 88.960 331.930 89.130 ;
        RECT 332.120 88.960 332.290 89.130 ;
        RECT 263.280 88.670 263.450 88.840 ;
        RECT 266.310 88.670 266.480 88.840 ;
        RECT 205.435 87.910 205.605 88.080 ;
        RECT 205.795 87.910 205.965 88.080 ;
        RECT 206.155 87.910 206.325 88.080 ;
        RECT 206.515 87.910 206.685 88.080 ;
        RECT 206.875 87.910 207.045 88.080 ;
        RECT 207.235 87.910 207.405 88.080 ;
        RECT 252.430 87.910 252.600 88.080 ;
        RECT 252.790 87.910 252.960 88.080 ;
        RECT 253.150 87.910 253.320 88.080 ;
        RECT 253.510 87.910 253.680 88.080 ;
        RECT 253.870 87.910 254.040 88.080 ;
        RECT 254.230 87.910 254.400 88.080 ;
        RECT 270.600 88.060 270.770 88.230 ;
        RECT 273.290 88.060 273.460 88.230 ;
        RECT 276.920 88.050 277.090 88.220 ;
        RECT 283.325 88.130 283.495 88.300 ;
        RECT 283.685 88.130 283.855 88.300 ;
        RECT 284.045 88.130 284.215 88.300 ;
        RECT 284.405 88.130 284.575 88.300 ;
        RECT 284.765 88.130 284.935 88.300 ;
        RECT 285.125 88.130 285.295 88.300 ;
        RECT 330.320 88.130 330.490 88.300 ;
        RECT 330.680 88.130 330.850 88.300 ;
        RECT 331.040 88.130 331.210 88.300 ;
        RECT 331.400 88.130 331.570 88.300 ;
        RECT 331.760 88.130 331.930 88.300 ;
        RECT 332.120 88.130 332.290 88.300 ;
        RECT 270.115 87.665 270.285 87.835 ;
        RECT 273.775 87.665 273.945 87.835 ;
        RECT 277.405 87.655 277.575 87.825 ;
        RECT 205.435 87.080 205.605 87.250 ;
        RECT 205.795 87.080 205.965 87.250 ;
        RECT 206.155 87.080 206.325 87.250 ;
        RECT 206.515 87.080 206.685 87.250 ;
        RECT 206.875 87.080 207.045 87.250 ;
        RECT 207.235 87.080 207.405 87.250 ;
        RECT 270.600 87.270 270.770 87.440 ;
        RECT 283.325 87.300 283.495 87.470 ;
        RECT 283.685 87.300 283.855 87.470 ;
        RECT 284.045 87.300 284.215 87.470 ;
        RECT 284.405 87.300 284.575 87.470 ;
        RECT 284.765 87.300 284.935 87.470 ;
        RECT 285.125 87.300 285.295 87.470 ;
        RECT 252.430 87.080 252.600 87.250 ;
        RECT 252.790 87.080 252.960 87.250 ;
        RECT 253.150 87.080 253.320 87.250 ;
        RECT 253.510 87.080 253.680 87.250 ;
        RECT 253.870 87.080 254.040 87.250 ;
        RECT 254.230 87.080 254.400 87.250 ;
        RECT 330.320 87.300 330.490 87.470 ;
        RECT 330.680 87.300 330.850 87.470 ;
        RECT 331.040 87.300 331.210 87.470 ;
        RECT 331.400 87.300 331.570 87.470 ;
        RECT 331.760 87.300 331.930 87.470 ;
        RECT 332.120 87.300 332.290 87.470 ;
        RECT 205.435 86.250 205.605 86.420 ;
        RECT 205.795 86.250 205.965 86.420 ;
        RECT 206.155 86.250 206.325 86.420 ;
        RECT 206.515 86.250 206.685 86.420 ;
        RECT 206.875 86.250 207.045 86.420 ;
        RECT 207.235 86.250 207.405 86.420 ;
        RECT 252.430 86.250 252.600 86.420 ;
        RECT 252.790 86.250 252.960 86.420 ;
        RECT 253.150 86.250 253.320 86.420 ;
        RECT 253.510 86.250 253.680 86.420 ;
        RECT 253.870 86.250 254.040 86.420 ;
        RECT 254.230 86.250 254.400 86.420 ;
        RECT 263.280 86.380 263.450 86.550 ;
        RECT 266.310 86.380 266.480 86.550 ;
        RECT 283.325 86.470 283.495 86.640 ;
        RECT 283.685 86.470 283.855 86.640 ;
        RECT 284.045 86.470 284.215 86.640 ;
        RECT 284.405 86.470 284.575 86.640 ;
        RECT 284.765 86.470 284.935 86.640 ;
        RECT 285.125 86.470 285.295 86.640 ;
        RECT 330.320 86.470 330.490 86.640 ;
        RECT 330.680 86.470 330.850 86.640 ;
        RECT 331.040 86.470 331.210 86.640 ;
        RECT 331.400 86.470 331.570 86.640 ;
        RECT 331.760 86.470 331.930 86.640 ;
        RECT 332.120 86.470 332.290 86.640 ;
        RECT 262.750 85.985 262.920 86.155 ;
        RECT 266.840 85.985 267.010 86.155 ;
        RECT 205.435 85.420 205.605 85.590 ;
        RECT 205.795 85.420 205.965 85.590 ;
        RECT 206.155 85.420 206.325 85.590 ;
        RECT 206.515 85.420 206.685 85.590 ;
        RECT 206.875 85.420 207.045 85.590 ;
        RECT 207.235 85.420 207.405 85.590 ;
        RECT 252.430 85.420 252.600 85.590 ;
        RECT 252.790 85.420 252.960 85.590 ;
        RECT 253.150 85.420 253.320 85.590 ;
        RECT 253.510 85.420 253.680 85.590 ;
        RECT 253.870 85.420 254.040 85.590 ;
        RECT 254.230 85.420 254.400 85.590 ;
        RECT 283.325 85.640 283.495 85.810 ;
        RECT 283.685 85.640 283.855 85.810 ;
        RECT 284.045 85.640 284.215 85.810 ;
        RECT 284.405 85.640 284.575 85.810 ;
        RECT 284.765 85.640 284.935 85.810 ;
        RECT 285.125 85.640 285.295 85.810 ;
        RECT 330.320 85.640 330.490 85.810 ;
        RECT 330.680 85.640 330.850 85.810 ;
        RECT 331.040 85.640 331.210 85.810 ;
        RECT 331.400 85.640 331.570 85.810 ;
        RECT 331.760 85.640 331.930 85.810 ;
        RECT 332.120 85.640 332.290 85.810 ;
        RECT 270.600 85.280 270.770 85.450 ;
        RECT 273.290 85.280 273.460 85.450 ;
        RECT 276.920 85.270 277.090 85.440 ;
        RECT 270.115 84.885 270.285 85.055 ;
        RECT 252.430 84.590 252.600 84.760 ;
        RECT 252.790 84.590 252.960 84.760 ;
        RECT 253.150 84.590 253.320 84.760 ;
        RECT 253.510 84.590 253.680 84.760 ;
        RECT 253.870 84.590 254.040 84.760 ;
        RECT 254.230 84.590 254.400 84.760 ;
        RECT 273.775 84.885 273.945 85.055 ;
        RECT 277.405 84.875 277.575 85.045 ;
        RECT 283.325 84.810 283.495 84.980 ;
        RECT 283.685 84.810 283.855 84.980 ;
        RECT 284.045 84.810 284.215 84.980 ;
        RECT 284.405 84.810 284.575 84.980 ;
        RECT 284.765 84.810 284.935 84.980 ;
        RECT 285.125 84.810 285.295 84.980 ;
        RECT 330.320 84.810 330.490 84.980 ;
        RECT 330.680 84.810 330.850 84.980 ;
        RECT 331.040 84.810 331.210 84.980 ;
        RECT 331.400 84.810 331.570 84.980 ;
        RECT 331.760 84.810 331.930 84.980 ;
        RECT 332.120 84.810 332.290 84.980 ;
        RECT 270.600 84.490 270.770 84.660 ;
        RECT 276.920 84.480 277.090 84.650 ;
        RECT 283.325 83.980 283.495 84.150 ;
        RECT 283.685 83.980 283.855 84.150 ;
        RECT 284.045 83.980 284.215 84.150 ;
        RECT 284.405 83.980 284.575 84.150 ;
        RECT 284.765 83.980 284.935 84.150 ;
        RECT 285.125 83.980 285.295 84.150 ;
        RECT 330.320 83.980 330.490 84.150 ;
        RECT 330.680 83.980 330.850 84.150 ;
        RECT 331.040 83.980 331.210 84.150 ;
        RECT 331.400 83.980 331.570 84.150 ;
        RECT 331.760 83.980 331.930 84.150 ;
        RECT 332.120 83.980 332.290 84.150 ;
        RECT 283.325 83.150 283.495 83.320 ;
        RECT 283.685 83.150 283.855 83.320 ;
        RECT 284.045 83.150 284.215 83.320 ;
        RECT 284.405 83.150 284.575 83.320 ;
        RECT 284.765 83.150 284.935 83.320 ;
        RECT 285.125 83.150 285.295 83.320 ;
        RECT 330.320 83.150 330.490 83.320 ;
        RECT 330.680 83.150 330.850 83.320 ;
        RECT 331.040 83.150 331.210 83.320 ;
        RECT 331.400 83.150 331.570 83.320 ;
        RECT 331.760 83.150 331.930 83.320 ;
        RECT 332.120 83.150 332.290 83.320 ;
        RECT 283.325 82.320 283.495 82.490 ;
        RECT 283.685 82.320 283.855 82.490 ;
        RECT 284.045 82.320 284.215 82.490 ;
        RECT 284.405 82.320 284.575 82.490 ;
        RECT 284.765 82.320 284.935 82.490 ;
        RECT 285.125 82.320 285.295 82.490 ;
        RECT 330.320 82.320 330.490 82.490 ;
        RECT 330.680 82.320 330.850 82.490 ;
        RECT 331.040 82.320 331.210 82.490 ;
        RECT 331.400 82.320 331.570 82.490 ;
        RECT 331.760 82.320 331.930 82.490 ;
        RECT 332.120 82.320 332.290 82.490 ;
        RECT 205.485 81.590 205.655 81.760 ;
        RECT 205.845 81.590 206.015 81.760 ;
        RECT 206.205 81.590 206.375 81.760 ;
        RECT 206.565 81.590 206.735 81.760 ;
        RECT 206.925 81.590 207.095 81.760 ;
        RECT 207.285 81.590 207.455 81.760 ;
        RECT 252.480 81.590 252.650 81.760 ;
        RECT 252.840 81.590 253.010 81.760 ;
        RECT 253.200 81.590 253.370 81.760 ;
        RECT 253.560 81.590 253.730 81.760 ;
        RECT 253.920 81.590 254.090 81.760 ;
        RECT 254.280 81.590 254.450 81.760 ;
        RECT 283.325 81.490 283.495 81.660 ;
        RECT 283.685 81.490 283.855 81.660 ;
        RECT 284.045 81.490 284.215 81.660 ;
        RECT 284.405 81.490 284.575 81.660 ;
        RECT 284.765 81.490 284.935 81.660 ;
        RECT 285.125 81.490 285.295 81.660 ;
        RECT 330.320 81.490 330.490 81.660 ;
        RECT 330.680 81.490 330.850 81.660 ;
        RECT 331.040 81.490 331.210 81.660 ;
        RECT 331.400 81.490 331.570 81.660 ;
        RECT 331.760 81.490 331.930 81.660 ;
        RECT 332.120 81.490 332.290 81.660 ;
        RECT 205.485 80.760 205.655 80.930 ;
        RECT 205.845 80.760 206.015 80.930 ;
        RECT 206.205 80.760 206.375 80.930 ;
        RECT 206.565 80.760 206.735 80.930 ;
        RECT 206.925 80.760 207.095 80.930 ;
        RECT 207.285 80.760 207.455 80.930 ;
        RECT 252.480 80.760 252.650 80.930 ;
        RECT 252.840 80.760 253.010 80.930 ;
        RECT 253.200 80.760 253.370 80.930 ;
        RECT 253.560 80.760 253.730 80.930 ;
        RECT 253.920 80.760 254.090 80.930 ;
        RECT 254.280 80.760 254.450 80.930 ;
        RECT 283.325 80.660 283.495 80.830 ;
        RECT 283.685 80.660 283.855 80.830 ;
        RECT 284.045 80.660 284.215 80.830 ;
        RECT 284.405 80.660 284.575 80.830 ;
        RECT 284.765 80.660 284.935 80.830 ;
        RECT 285.125 80.660 285.295 80.830 ;
        RECT 330.320 80.660 330.490 80.830 ;
        RECT 330.680 80.660 330.850 80.830 ;
        RECT 331.040 80.660 331.210 80.830 ;
        RECT 331.400 80.660 331.570 80.830 ;
        RECT 331.760 80.660 331.930 80.830 ;
        RECT 332.120 80.660 332.290 80.830 ;
        RECT 205.485 79.930 205.655 80.100 ;
        RECT 205.845 79.930 206.015 80.100 ;
        RECT 206.205 79.930 206.375 80.100 ;
        RECT 206.565 79.930 206.735 80.100 ;
        RECT 206.925 79.930 207.095 80.100 ;
        RECT 207.285 79.930 207.455 80.100 ;
        RECT 252.480 79.930 252.650 80.100 ;
        RECT 252.840 79.930 253.010 80.100 ;
        RECT 253.200 79.930 253.370 80.100 ;
        RECT 253.560 79.930 253.730 80.100 ;
        RECT 253.920 79.930 254.090 80.100 ;
        RECT 254.280 79.930 254.450 80.100 ;
        RECT 205.485 79.100 205.655 79.270 ;
        RECT 205.845 79.100 206.015 79.270 ;
        RECT 206.205 79.100 206.375 79.270 ;
        RECT 206.565 79.100 206.735 79.270 ;
        RECT 206.925 79.100 207.095 79.270 ;
        RECT 207.285 79.100 207.455 79.270 ;
        RECT 252.480 79.100 252.650 79.270 ;
        RECT 252.840 79.100 253.010 79.270 ;
        RECT 253.200 79.100 253.370 79.270 ;
        RECT 253.560 79.100 253.730 79.270 ;
        RECT 253.920 79.100 254.090 79.270 ;
        RECT 254.280 79.100 254.450 79.270 ;
        RECT 205.485 78.270 205.655 78.440 ;
        RECT 205.845 78.270 206.015 78.440 ;
        RECT 206.205 78.270 206.375 78.440 ;
        RECT 206.565 78.270 206.735 78.440 ;
        RECT 206.925 78.270 207.095 78.440 ;
        RECT 207.285 78.270 207.455 78.440 ;
        RECT 252.480 78.270 252.650 78.440 ;
        RECT 252.840 78.270 253.010 78.440 ;
        RECT 253.200 78.270 253.370 78.440 ;
        RECT 253.560 78.270 253.730 78.440 ;
        RECT 253.920 78.270 254.090 78.440 ;
        RECT 254.280 78.270 254.450 78.440 ;
        RECT 205.485 77.440 205.655 77.610 ;
        RECT 205.845 77.440 206.015 77.610 ;
        RECT 206.205 77.440 206.375 77.610 ;
        RECT 206.565 77.440 206.735 77.610 ;
        RECT 206.925 77.440 207.095 77.610 ;
        RECT 207.285 77.440 207.455 77.610 ;
        RECT 252.480 77.440 252.650 77.610 ;
        RECT 252.840 77.440 253.010 77.610 ;
        RECT 253.200 77.440 253.370 77.610 ;
        RECT 253.560 77.440 253.730 77.610 ;
        RECT 253.920 77.440 254.090 77.610 ;
        RECT 254.280 77.440 254.450 77.610 ;
        RECT 205.485 76.610 205.655 76.780 ;
        RECT 205.845 76.610 206.015 76.780 ;
        RECT 206.205 76.610 206.375 76.780 ;
        RECT 206.565 76.610 206.735 76.780 ;
        RECT 206.925 76.610 207.095 76.780 ;
        RECT 207.285 76.610 207.455 76.780 ;
        RECT 252.480 76.610 252.650 76.780 ;
        RECT 252.840 76.610 253.010 76.780 ;
        RECT 253.200 76.610 253.370 76.780 ;
        RECT 253.560 76.610 253.730 76.780 ;
        RECT 253.920 76.610 254.090 76.780 ;
        RECT 254.280 76.610 254.450 76.780 ;
        RECT 205.485 75.780 205.655 75.950 ;
        RECT 205.845 75.780 206.015 75.950 ;
        RECT 206.205 75.780 206.375 75.950 ;
        RECT 206.565 75.780 206.735 75.950 ;
        RECT 206.925 75.780 207.095 75.950 ;
        RECT 207.285 75.780 207.455 75.950 ;
        RECT 252.480 75.780 252.650 75.950 ;
        RECT 252.840 75.780 253.010 75.950 ;
        RECT 253.200 75.780 253.370 75.950 ;
        RECT 253.560 75.780 253.730 75.950 ;
        RECT 253.920 75.780 254.090 75.950 ;
        RECT 254.280 75.780 254.450 75.950 ;
        RECT 205.485 74.950 205.655 75.120 ;
        RECT 205.845 74.950 206.015 75.120 ;
        RECT 206.205 74.950 206.375 75.120 ;
        RECT 206.565 74.950 206.735 75.120 ;
        RECT 206.925 74.950 207.095 75.120 ;
        RECT 207.285 74.950 207.455 75.120 ;
        RECT 252.480 74.950 252.650 75.120 ;
        RECT 252.840 74.950 253.010 75.120 ;
        RECT 253.200 74.950 253.370 75.120 ;
        RECT 253.560 74.950 253.730 75.120 ;
        RECT 253.920 74.950 254.090 75.120 ;
        RECT 254.280 74.950 254.450 75.120 ;
        RECT 263.330 79.100 263.500 79.270 ;
        RECT 266.680 79.100 266.850 79.270 ;
        RECT 271.190 79.100 271.360 79.270 ;
        RECT 274.540 79.100 274.710 79.270 ;
        RECT 259.350 78.695 259.520 78.865 ;
        RECT 260.320 78.695 260.490 78.865 ;
        RECT 262.800 78.705 262.970 78.875 ;
        RECT 263.860 78.705 264.030 78.875 ;
        RECT 266.150 78.705 266.320 78.875 ;
        RECT 267.210 78.705 267.380 78.875 ;
        RECT 270.660 78.705 270.830 78.875 ;
        RECT 271.720 78.705 271.890 78.875 ;
        RECT 274.010 78.705 274.180 78.875 ;
        RECT 275.070 78.705 275.240 78.875 ;
        RECT 277.550 78.695 277.720 78.865 ;
        RECT 278.520 78.695 278.690 78.865 ;
        RECT 259.835 78.300 260.005 78.470 ;
        RECT 263.330 78.310 263.500 78.480 ;
        RECT 274.540 78.310 274.710 78.480 ;
        RECT 278.035 78.300 278.205 78.470 ;
        RECT 259.825 76.060 259.995 76.230 ;
        RECT 263.340 76.050 263.510 76.220 ;
        RECT 274.530 76.050 274.700 76.220 ;
        RECT 278.045 76.060 278.215 76.230 ;
        RECT 262.810 75.655 262.980 75.825 ;
        RECT 263.870 75.655 264.040 75.825 ;
        RECT 266.150 75.625 266.320 75.795 ;
        RECT 267.210 75.625 267.380 75.795 ;
        RECT 270.660 75.625 270.830 75.795 ;
        RECT 271.720 75.625 271.890 75.795 ;
        RECT 274.000 75.655 274.170 75.825 ;
        RECT 275.060 75.655 275.230 75.825 ;
        RECT 263.340 75.260 263.510 75.430 ;
        RECT 266.680 75.230 266.850 75.400 ;
        RECT 271.190 75.230 271.360 75.400 ;
        RECT 274.530 75.260 274.700 75.430 ;
        RECT 283.325 79.830 283.495 80.000 ;
        RECT 283.685 79.830 283.855 80.000 ;
        RECT 284.045 79.830 284.215 80.000 ;
        RECT 284.405 79.830 284.575 80.000 ;
        RECT 284.765 79.830 284.935 80.000 ;
        RECT 285.125 79.830 285.295 80.000 ;
        RECT 330.320 79.830 330.490 80.000 ;
        RECT 330.680 79.830 330.850 80.000 ;
        RECT 331.040 79.830 331.210 80.000 ;
        RECT 331.400 79.830 331.570 80.000 ;
        RECT 331.760 79.830 331.930 80.000 ;
        RECT 332.120 79.830 332.290 80.000 ;
        RECT 283.325 79.000 283.495 79.170 ;
        RECT 283.685 79.000 283.855 79.170 ;
        RECT 284.045 79.000 284.215 79.170 ;
        RECT 284.405 79.000 284.575 79.170 ;
        RECT 284.765 79.000 284.935 79.170 ;
        RECT 285.125 79.000 285.295 79.170 ;
        RECT 330.320 79.000 330.490 79.170 ;
        RECT 330.680 79.000 330.850 79.170 ;
        RECT 331.040 79.000 331.210 79.170 ;
        RECT 331.400 79.000 331.570 79.170 ;
        RECT 331.760 79.000 331.930 79.170 ;
        RECT 332.120 79.000 332.290 79.170 ;
        RECT 283.325 78.170 283.495 78.340 ;
        RECT 283.685 78.170 283.855 78.340 ;
        RECT 284.045 78.170 284.215 78.340 ;
        RECT 284.405 78.170 284.575 78.340 ;
        RECT 284.765 78.170 284.935 78.340 ;
        RECT 285.125 78.170 285.295 78.340 ;
        RECT 330.320 78.170 330.490 78.340 ;
        RECT 330.680 78.170 330.850 78.340 ;
        RECT 331.040 78.170 331.210 78.340 ;
        RECT 331.400 78.170 331.570 78.340 ;
        RECT 331.760 78.170 331.930 78.340 ;
        RECT 332.120 78.170 332.290 78.340 ;
        RECT 283.325 77.340 283.495 77.510 ;
        RECT 283.685 77.340 283.855 77.510 ;
        RECT 284.045 77.340 284.215 77.510 ;
        RECT 284.405 77.340 284.575 77.510 ;
        RECT 284.765 77.340 284.935 77.510 ;
        RECT 285.125 77.340 285.295 77.510 ;
        RECT 330.320 77.340 330.490 77.510 ;
        RECT 330.680 77.340 330.850 77.510 ;
        RECT 331.040 77.340 331.210 77.510 ;
        RECT 331.400 77.340 331.570 77.510 ;
        RECT 331.760 77.340 331.930 77.510 ;
        RECT 332.120 77.340 332.290 77.510 ;
        RECT 283.325 76.510 283.495 76.680 ;
        RECT 283.685 76.510 283.855 76.680 ;
        RECT 284.045 76.510 284.215 76.680 ;
        RECT 284.405 76.510 284.575 76.680 ;
        RECT 284.765 76.510 284.935 76.680 ;
        RECT 285.125 76.510 285.295 76.680 ;
        RECT 330.320 76.510 330.490 76.680 ;
        RECT 330.680 76.510 330.850 76.680 ;
        RECT 331.040 76.510 331.210 76.680 ;
        RECT 331.400 76.510 331.570 76.680 ;
        RECT 331.760 76.510 331.930 76.680 ;
        RECT 332.120 76.510 332.290 76.680 ;
        RECT 283.325 75.680 283.495 75.850 ;
        RECT 283.685 75.680 283.855 75.850 ;
        RECT 284.045 75.680 284.215 75.850 ;
        RECT 284.405 75.680 284.575 75.850 ;
        RECT 284.765 75.680 284.935 75.850 ;
        RECT 285.125 75.680 285.295 75.850 ;
        RECT 330.320 75.680 330.490 75.850 ;
        RECT 330.680 75.680 330.850 75.850 ;
        RECT 331.040 75.680 331.210 75.850 ;
        RECT 331.400 75.680 331.570 75.850 ;
        RECT 331.760 75.680 331.930 75.850 ;
        RECT 332.120 75.680 332.290 75.850 ;
        RECT 283.325 74.850 283.495 75.020 ;
        RECT 283.685 74.850 283.855 75.020 ;
        RECT 284.045 74.850 284.215 75.020 ;
        RECT 284.405 74.850 284.575 75.020 ;
        RECT 284.765 74.850 284.935 75.020 ;
        RECT 285.125 74.850 285.295 75.020 ;
        RECT 330.320 74.850 330.490 75.020 ;
        RECT 330.680 74.850 330.850 75.020 ;
        RECT 331.040 74.850 331.210 75.020 ;
        RECT 331.400 74.850 331.570 75.020 ;
        RECT 331.760 74.850 331.930 75.020 ;
        RECT 332.120 74.850 332.290 75.020 ;
        RECT 205.485 74.120 205.655 74.290 ;
        RECT 205.845 74.120 206.015 74.290 ;
        RECT 206.205 74.120 206.375 74.290 ;
        RECT 206.565 74.120 206.735 74.290 ;
        RECT 206.925 74.120 207.095 74.290 ;
        RECT 207.285 74.120 207.455 74.290 ;
        RECT 252.480 74.120 252.650 74.290 ;
        RECT 252.840 74.120 253.010 74.290 ;
        RECT 253.200 74.120 253.370 74.290 ;
        RECT 253.560 74.120 253.730 74.290 ;
        RECT 253.920 74.120 254.090 74.290 ;
        RECT 254.280 74.120 254.450 74.290 ;
        RECT 283.325 74.020 283.495 74.190 ;
        RECT 283.685 74.020 283.855 74.190 ;
        RECT 284.045 74.020 284.215 74.190 ;
        RECT 284.405 74.020 284.575 74.190 ;
        RECT 284.765 74.020 284.935 74.190 ;
        RECT 285.125 74.020 285.295 74.190 ;
        RECT 330.320 74.020 330.490 74.190 ;
        RECT 330.680 74.020 330.850 74.190 ;
        RECT 331.040 74.020 331.210 74.190 ;
        RECT 331.400 74.020 331.570 74.190 ;
        RECT 331.760 74.020 331.930 74.190 ;
        RECT 332.120 74.020 332.290 74.190 ;
        RECT 205.485 73.290 205.655 73.460 ;
        RECT 205.845 73.290 206.015 73.460 ;
        RECT 206.205 73.290 206.375 73.460 ;
        RECT 206.565 73.290 206.735 73.460 ;
        RECT 206.925 73.290 207.095 73.460 ;
        RECT 207.285 73.290 207.455 73.460 ;
        RECT 252.480 73.290 252.650 73.460 ;
        RECT 252.840 73.290 253.010 73.460 ;
        RECT 253.200 73.290 253.370 73.460 ;
        RECT 253.560 73.290 253.730 73.460 ;
        RECT 253.920 73.290 254.090 73.460 ;
        RECT 254.280 73.290 254.450 73.460 ;
        RECT 283.325 73.190 283.495 73.360 ;
        RECT 283.685 73.190 283.855 73.360 ;
        RECT 284.045 73.190 284.215 73.360 ;
        RECT 284.405 73.190 284.575 73.360 ;
        RECT 284.765 73.190 284.935 73.360 ;
        RECT 285.125 73.190 285.295 73.360 ;
        RECT 330.320 73.190 330.490 73.360 ;
        RECT 330.680 73.190 330.850 73.360 ;
        RECT 331.040 73.190 331.210 73.360 ;
        RECT 331.400 73.190 331.570 73.360 ;
        RECT 331.760 73.190 331.930 73.360 ;
        RECT 332.120 73.190 332.290 73.360 ;
        RECT 205.485 72.460 205.655 72.630 ;
        RECT 205.845 72.460 206.015 72.630 ;
        RECT 206.205 72.460 206.375 72.630 ;
        RECT 206.565 72.460 206.735 72.630 ;
        RECT 206.925 72.460 207.095 72.630 ;
        RECT 207.285 72.460 207.455 72.630 ;
        RECT 252.480 72.460 252.650 72.630 ;
        RECT 252.840 72.460 253.010 72.630 ;
        RECT 253.200 72.460 253.370 72.630 ;
        RECT 253.560 72.460 253.730 72.630 ;
        RECT 253.920 72.460 254.090 72.630 ;
        RECT 254.280 72.460 254.450 72.630 ;
        RECT 283.325 72.360 283.495 72.530 ;
        RECT 283.685 72.360 283.855 72.530 ;
        RECT 284.045 72.360 284.215 72.530 ;
        RECT 284.405 72.360 284.575 72.530 ;
        RECT 284.765 72.360 284.935 72.530 ;
        RECT 285.125 72.360 285.295 72.530 ;
        RECT 330.320 72.360 330.490 72.530 ;
        RECT 330.680 72.360 330.850 72.530 ;
        RECT 331.040 72.360 331.210 72.530 ;
        RECT 331.400 72.360 331.570 72.530 ;
        RECT 331.760 72.360 331.930 72.530 ;
        RECT 332.120 72.360 332.290 72.530 ;
        RECT 205.485 71.630 205.655 71.800 ;
        RECT 205.845 71.630 206.015 71.800 ;
        RECT 206.205 71.630 206.375 71.800 ;
        RECT 206.565 71.630 206.735 71.800 ;
        RECT 206.925 71.630 207.095 71.800 ;
        RECT 207.285 71.630 207.455 71.800 ;
        RECT 252.480 71.630 252.650 71.800 ;
        RECT 252.840 71.630 253.010 71.800 ;
        RECT 253.200 71.630 253.370 71.800 ;
        RECT 253.560 71.630 253.730 71.800 ;
        RECT 253.920 71.630 254.090 71.800 ;
        RECT 254.280 71.630 254.450 71.800 ;
        RECT 283.325 71.530 283.495 71.700 ;
        RECT 283.685 71.530 283.855 71.700 ;
        RECT 284.045 71.530 284.215 71.700 ;
        RECT 284.405 71.530 284.575 71.700 ;
        RECT 284.765 71.530 284.935 71.700 ;
        RECT 285.125 71.530 285.295 71.700 ;
        RECT 330.320 71.530 330.490 71.700 ;
        RECT 330.680 71.530 330.850 71.700 ;
        RECT 331.040 71.530 331.210 71.700 ;
        RECT 331.400 71.530 331.570 71.700 ;
        RECT 331.760 71.530 331.930 71.700 ;
        RECT 332.120 71.530 332.290 71.700 ;
        RECT 205.485 70.800 205.655 70.970 ;
        RECT 205.845 70.800 206.015 70.970 ;
        RECT 206.205 70.800 206.375 70.970 ;
        RECT 206.565 70.800 206.735 70.970 ;
        RECT 206.925 70.800 207.095 70.970 ;
        RECT 207.285 70.800 207.455 70.970 ;
        RECT 252.480 70.800 252.650 70.970 ;
        RECT 252.840 70.800 253.010 70.970 ;
        RECT 253.200 70.800 253.370 70.970 ;
        RECT 253.560 70.800 253.730 70.970 ;
        RECT 253.920 70.800 254.090 70.970 ;
        RECT 254.280 70.800 254.450 70.970 ;
        RECT 274.115 70.400 276.085 70.930 ;
        RECT 283.325 70.700 283.495 70.870 ;
        RECT 283.685 70.700 283.855 70.870 ;
        RECT 284.045 70.700 284.215 70.870 ;
        RECT 284.405 70.700 284.575 70.870 ;
        RECT 284.765 70.700 284.935 70.870 ;
        RECT 285.125 70.700 285.295 70.870 ;
        RECT 330.320 70.700 330.490 70.870 ;
        RECT 330.680 70.700 330.850 70.870 ;
        RECT 331.040 70.700 331.210 70.870 ;
        RECT 331.400 70.700 331.570 70.870 ;
        RECT 331.760 70.700 331.930 70.870 ;
        RECT 332.120 70.700 332.290 70.870 ;
        RECT 205.485 69.970 205.655 70.140 ;
        RECT 205.845 69.970 206.015 70.140 ;
        RECT 206.205 69.970 206.375 70.140 ;
        RECT 206.565 69.970 206.735 70.140 ;
        RECT 206.925 69.970 207.095 70.140 ;
        RECT 207.285 69.970 207.455 70.140 ;
        RECT 252.480 69.970 252.650 70.140 ;
        RECT 252.840 69.970 253.010 70.140 ;
        RECT 253.200 69.970 253.370 70.140 ;
        RECT 253.560 69.970 253.730 70.140 ;
        RECT 253.920 69.970 254.090 70.140 ;
        RECT 254.280 69.970 254.450 70.140 ;
        RECT 283.325 69.870 283.495 70.040 ;
        RECT 283.685 69.870 283.855 70.040 ;
        RECT 284.045 69.870 284.215 70.040 ;
        RECT 284.405 69.870 284.575 70.040 ;
        RECT 284.765 69.870 284.935 70.040 ;
        RECT 285.125 69.870 285.295 70.040 ;
        RECT 330.320 69.870 330.490 70.040 ;
        RECT 330.680 69.870 330.850 70.040 ;
        RECT 331.040 69.870 331.210 70.040 ;
        RECT 331.400 69.870 331.570 70.040 ;
        RECT 331.760 69.870 331.930 70.040 ;
        RECT 332.120 69.870 332.290 70.040 ;
        RECT 205.485 69.140 205.655 69.310 ;
        RECT 205.845 69.140 206.015 69.310 ;
        RECT 206.205 69.140 206.375 69.310 ;
        RECT 206.565 69.140 206.735 69.310 ;
        RECT 206.925 69.140 207.095 69.310 ;
        RECT 207.285 69.140 207.455 69.310 ;
        RECT 252.480 69.140 252.650 69.310 ;
        RECT 252.840 69.140 253.010 69.310 ;
        RECT 253.200 69.140 253.370 69.310 ;
        RECT 253.560 69.140 253.730 69.310 ;
        RECT 253.920 69.140 254.090 69.310 ;
        RECT 254.280 69.140 254.450 69.310 ;
        RECT 283.325 69.040 283.495 69.210 ;
        RECT 283.685 69.040 283.855 69.210 ;
        RECT 284.045 69.040 284.215 69.210 ;
        RECT 284.405 69.040 284.575 69.210 ;
        RECT 284.765 69.040 284.935 69.210 ;
        RECT 285.125 69.040 285.295 69.210 ;
        RECT 330.320 69.040 330.490 69.210 ;
        RECT 330.680 69.040 330.850 69.210 ;
        RECT 331.040 69.040 331.210 69.210 ;
        RECT 331.400 69.040 331.570 69.210 ;
        RECT 331.760 69.040 331.930 69.210 ;
        RECT 332.120 69.040 332.290 69.210 ;
        RECT 205.485 68.310 205.655 68.480 ;
        RECT 205.845 68.310 206.015 68.480 ;
        RECT 206.205 68.310 206.375 68.480 ;
        RECT 206.565 68.310 206.735 68.480 ;
        RECT 206.925 68.310 207.095 68.480 ;
        RECT 207.285 68.310 207.455 68.480 ;
        RECT 252.480 68.310 252.650 68.480 ;
        RECT 252.840 68.310 253.010 68.480 ;
        RECT 253.200 68.310 253.370 68.480 ;
        RECT 253.560 68.310 253.730 68.480 ;
        RECT 253.920 68.310 254.090 68.480 ;
        RECT 254.280 68.310 254.450 68.480 ;
        RECT 283.325 68.210 283.495 68.380 ;
        RECT 283.685 68.210 283.855 68.380 ;
        RECT 284.045 68.210 284.215 68.380 ;
        RECT 284.405 68.210 284.575 68.380 ;
        RECT 284.765 68.210 284.935 68.380 ;
        RECT 285.125 68.210 285.295 68.380 ;
        RECT 330.320 68.210 330.490 68.380 ;
        RECT 330.680 68.210 330.850 68.380 ;
        RECT 331.040 68.210 331.210 68.380 ;
        RECT 331.400 68.210 331.570 68.380 ;
        RECT 331.760 68.210 331.930 68.380 ;
        RECT 332.120 68.210 332.290 68.380 ;
        RECT 205.485 67.480 205.655 67.650 ;
        RECT 205.845 67.480 206.015 67.650 ;
        RECT 206.205 67.480 206.375 67.650 ;
        RECT 206.565 67.480 206.735 67.650 ;
        RECT 206.925 67.480 207.095 67.650 ;
        RECT 207.285 67.480 207.455 67.650 ;
        RECT 252.480 67.480 252.650 67.650 ;
        RECT 252.840 67.480 253.010 67.650 ;
        RECT 253.200 67.480 253.370 67.650 ;
        RECT 253.560 67.480 253.730 67.650 ;
        RECT 253.920 67.480 254.090 67.650 ;
        RECT 254.280 67.480 254.450 67.650 ;
        RECT 261.265 67.610 261.435 67.780 ;
        RECT 261.625 67.610 261.795 67.780 ;
        RECT 264.455 67.610 264.625 67.780 ;
        RECT 264.815 67.610 264.985 67.780 ;
        RECT 273.055 67.610 273.225 67.780 ;
        RECT 273.415 67.610 273.585 67.780 ;
        RECT 276.245 67.610 276.415 67.780 ;
        RECT 276.605 67.610 276.775 67.780 ;
        RECT 283.325 67.380 283.495 67.550 ;
        RECT 283.685 67.380 283.855 67.550 ;
        RECT 284.045 67.380 284.215 67.550 ;
        RECT 284.405 67.380 284.575 67.550 ;
        RECT 284.765 67.380 284.935 67.550 ;
        RECT 285.125 67.380 285.295 67.550 ;
        RECT 330.320 67.380 330.490 67.550 ;
        RECT 330.680 67.380 330.850 67.550 ;
        RECT 331.040 67.380 331.210 67.550 ;
        RECT 331.400 67.380 331.570 67.550 ;
        RECT 331.760 67.380 331.930 67.550 ;
        RECT 332.120 67.380 332.290 67.550 ;
        RECT 267.885 66.965 268.055 67.135 ;
        RECT 252.480 66.650 252.650 66.820 ;
        RECT 252.840 66.650 253.010 66.820 ;
        RECT 253.200 66.650 253.370 66.820 ;
        RECT 253.560 66.650 253.730 66.820 ;
        RECT 253.920 66.650 254.090 66.820 ;
        RECT 254.280 66.650 254.450 66.820 ;
        RECT 268.410 66.745 268.580 66.915 ;
        RECT 283.325 66.550 283.495 66.720 ;
        RECT 283.685 66.550 283.855 66.720 ;
        RECT 284.045 66.550 284.215 66.720 ;
        RECT 284.405 66.550 284.575 66.720 ;
        RECT 284.765 66.550 284.935 66.720 ;
        RECT 285.125 66.550 285.295 66.720 ;
        RECT 330.320 66.550 330.490 66.720 ;
        RECT 330.680 66.550 330.850 66.720 ;
        RECT 331.040 66.550 331.210 66.720 ;
        RECT 331.400 66.550 331.570 66.720 ;
        RECT 331.760 66.550 331.930 66.720 ;
        RECT 332.120 66.550 332.290 66.720 ;
        RECT 268.410 65.120 268.580 65.290 ;
        RECT 265.140 64.900 265.310 65.070 ;
        RECT 264.140 64.680 264.310 64.850 ;
        RECT 264.500 64.680 264.670 64.850 ;
        RECT 270.175 64.900 270.345 65.070 ;
        RECT 268.410 64.680 268.580 64.850 ;
        RECT 270.660 64.680 270.830 64.850 ;
      LAYER met1 ;
        RECT 279.250 133.100 280.250 134.100 ;
        RECT 205.335 130.150 207.495 131.330 ;
        RECT 252.335 130.980 256.165 131.330 ;
        RECT 205.335 128.490 207.495 129.670 ;
        RECT 252.335 129.320 254.495 130.500 ;
        RECT 205.335 126.830 207.495 128.010 ;
        RECT 252.335 127.660 254.495 128.840 ;
        RECT 205.335 125.170 207.495 126.350 ;
        RECT 252.335 126.000 254.495 127.180 ;
        RECT 205.335 123.510 207.495 124.690 ;
        RECT 252.335 124.340 254.495 125.520 ;
        RECT 205.335 121.850 207.495 123.030 ;
        RECT 252.335 122.680 254.495 123.860 ;
        RECT 205.335 120.190 207.495 121.370 ;
        RECT 252.335 121.020 254.495 122.200 ;
        RECT 205.335 118.530 207.495 119.710 ;
        RECT 252.335 119.360 254.495 120.540 ;
        RECT 205.335 116.870 207.495 118.050 ;
        RECT 252.335 117.700 254.495 118.880 ;
        RECT 205.335 115.210 207.495 116.390 ;
        RECT 252.335 116.040 254.495 117.220 ;
        RECT 205.335 113.550 207.495 114.730 ;
        RECT 252.335 114.380 254.495 115.560 ;
        RECT 205.335 111.890 207.495 113.070 ;
        RECT 252.335 112.720 254.495 113.900 ;
        RECT 205.335 110.230 207.495 111.410 ;
        RECT 252.335 111.060 254.495 112.240 ;
        RECT 205.335 108.570 207.495 109.750 ;
        RECT 252.335 109.400 254.495 110.580 ;
        RECT 205.335 106.910 207.495 108.090 ;
        RECT 252.335 107.740 254.495 108.920 ;
        RECT 205.335 105.250 207.495 106.430 ;
        RECT 252.335 106.080 254.495 107.260 ;
        RECT 205.335 103.590 207.495 104.770 ;
        RECT 252.335 104.420 254.495 105.600 ;
        RECT 205.335 101.930 207.495 103.110 ;
        RECT 252.335 102.760 254.495 103.940 ;
        RECT 205.335 100.270 207.495 101.450 ;
        RECT 252.335 101.100 254.495 102.280 ;
        RECT 255.670 102.165 256.165 130.980 ;
        RECT 257.395 128.890 259.555 130.750 ;
        RECT 279.465 130.700 280.000 133.100 ;
        RECT 278.420 130.110 280.525 130.700 ;
        RECT 283.225 130.365 285.385 131.550 ;
        RECT 257.395 126.550 259.555 128.410 ;
        RECT 278.395 127.720 280.555 129.580 ;
        RECT 283.225 128.710 285.385 129.895 ;
        RECT 330.225 129.540 332.385 130.720 ;
        RECT 257.395 124.210 259.555 126.070 ;
        RECT 278.395 125.380 280.555 127.240 ;
        RECT 283.225 127.055 285.385 128.240 ;
        RECT 330.225 127.880 332.385 129.060 ;
        RECT 283.225 125.400 285.385 126.585 ;
        RECT 330.225 126.220 332.385 127.400 ;
        RECT 257.395 121.870 259.555 123.730 ;
        RECT 278.395 123.040 280.555 124.900 ;
        RECT 283.225 123.745 285.385 124.930 ;
        RECT 330.225 124.560 332.385 125.740 ;
        RECT 257.395 119.530 259.555 121.390 ;
        RECT 278.395 120.700 280.555 122.560 ;
        RECT 283.225 122.090 285.385 123.275 ;
        RECT 330.225 122.900 332.385 124.080 ;
        RECT 283.225 120.435 285.385 121.620 ;
        RECT 330.225 121.240 332.385 122.420 ;
        RECT 257.395 117.190 259.555 119.050 ;
        RECT 278.395 118.360 280.555 120.220 ;
        RECT 283.225 118.780 285.385 119.965 ;
        RECT 330.225 119.580 332.385 120.760 ;
        RECT 257.395 114.850 259.555 116.710 ;
        RECT 278.395 116.020 280.555 117.880 ;
        RECT 283.225 117.125 285.385 118.310 ;
        RECT 330.225 117.920 332.385 119.100 ;
        RECT 257.395 112.510 259.555 114.370 ;
        RECT 278.395 113.680 280.555 115.540 ;
        RECT 283.225 115.470 285.385 116.655 ;
        RECT 330.225 116.260 332.385 117.440 ;
        RECT 283.225 113.815 285.385 115.000 ;
        RECT 330.225 114.600 332.385 115.780 ;
        RECT 257.395 110.170 259.555 112.030 ;
        RECT 278.395 111.340 280.555 113.200 ;
        RECT 283.225 112.160 285.385 113.345 ;
        RECT 330.225 112.940 332.385 114.120 ;
        RECT 257.395 107.830 259.555 109.690 ;
        RECT 278.395 109.000 280.555 110.860 ;
        RECT 283.225 110.505 285.385 111.690 ;
        RECT 330.225 111.280 332.385 112.460 ;
        RECT 283.255 110.500 285.360 110.505 ;
        RECT 283.225 108.850 285.385 110.035 ;
        RECT 330.225 109.620 332.385 110.800 ;
        RECT 283.255 108.840 285.360 108.850 ;
        RECT 257.395 105.490 259.555 107.350 ;
        RECT 278.395 106.660 280.555 108.520 ;
        RECT 283.225 107.195 285.385 108.380 ;
        RECT 330.225 107.960 332.385 109.140 ;
        RECT 283.255 107.180 285.360 107.195 ;
        RECT 257.395 103.150 259.555 105.010 ;
        RECT 278.395 104.320 280.555 106.180 ;
        RECT 283.225 105.540 285.385 106.725 ;
        RECT 330.225 106.300 332.385 107.480 ;
        RECT 283.255 105.520 285.360 105.540 ;
        RECT 283.225 103.885 285.385 105.070 ;
        RECT 330.225 104.640 332.385 105.820 ;
        RECT 283.255 103.860 285.360 103.885 ;
        RECT 278.420 103.200 280.525 103.790 ;
        RECT 279.225 102.165 279.835 103.200 ;
        RECT 283.225 102.230 285.385 103.415 ;
        RECT 330.225 102.980 332.385 104.160 ;
        RECT 283.255 102.200 285.360 102.230 ;
        RECT 255.670 101.680 279.835 102.165 ;
        RECT 205.335 98.610 207.495 99.790 ;
        RECT 252.335 99.440 254.495 100.620 ;
        RECT 205.335 96.950 207.495 98.130 ;
        RECT 252.335 97.780 254.495 98.960 ;
        RECT 205.335 95.290 207.495 96.470 ;
        RECT 252.335 96.120 254.495 97.300 ;
        RECT 264.940 96.770 265.160 101.680 ;
        RECT 268.665 100.790 269.455 100.870 ;
        RECT 268.665 100.545 274.110 100.790 ;
        RECT 268.665 100.475 269.455 100.545 ;
        RECT 267.215 99.545 268.135 99.640 ;
        RECT 267.215 99.495 270.915 99.545 ;
        RECT 266.285 99.330 270.915 99.495 ;
        RECT 266.285 99.275 268.165 99.330 ;
        RECT 266.285 98.900 266.505 99.275 ;
        RECT 267.215 99.215 268.135 99.275 ;
        RECT 270.475 99.150 270.895 99.330 ;
        RECT 271.065 99.305 273.600 99.555 ;
        RECT 270.070 99.100 270.275 99.105 ;
        RECT 268.205 98.950 268.995 98.995 ;
        RECT 266.185 98.670 266.605 98.900 ;
        RECT 266.835 98.745 269.025 98.950 ;
        RECT 266.835 98.620 267.040 98.745 ;
        RECT 266.810 98.160 267.040 98.620 ;
        RECT 268.205 98.600 268.995 98.745 ;
        RECT 270.070 98.640 270.315 99.100 ;
        RECT 266.835 98.135 267.040 98.160 ;
        RECT 270.070 97.695 270.275 98.640 ;
        RECT 270.475 98.455 270.895 98.590 ;
        RECT 271.065 98.455 271.315 99.305 ;
        RECT 273.165 99.150 273.585 99.305 ;
        RECT 273.865 99.100 274.110 100.545 ;
        RECT 273.745 98.670 274.110 99.100 ;
        RECT 273.745 98.640 273.975 98.670 ;
        RECT 270.470 98.205 271.315 98.455 ;
        RECT 270.070 97.400 271.015 97.695 ;
        RECT 270.180 97.310 271.015 97.400 ;
        RECT 264.930 96.600 270.875 96.770 ;
        RECT 264.930 96.550 270.895 96.600 ;
        RECT 266.280 95.820 266.500 96.550 ;
        RECT 270.475 96.370 270.895 96.550 ;
        RECT 271.065 96.555 273.600 96.805 ;
        RECT 268.175 96.165 268.465 96.205 ;
        RECT 270.085 96.165 270.315 96.320 ;
        RECT 268.175 95.960 270.315 96.165 ;
        RECT 205.335 93.630 207.495 94.810 ;
        RECT 252.335 94.460 254.495 95.640 ;
        RECT 266.185 95.590 266.605 95.820 ;
        RECT 262.635 95.540 262.895 95.570 ;
        RECT 262.635 95.080 262.950 95.540 ;
        RECT 266.810 95.430 267.040 95.540 ;
        RECT 268.175 95.430 268.465 95.960 ;
        RECT 270.085 95.860 270.315 95.960 ;
        RECT 270.475 95.680 270.895 95.810 ;
        RECT 271.065 95.680 271.315 96.555 ;
        RECT 273.165 96.370 273.585 96.555 ;
        RECT 273.880 96.320 274.170 96.330 ;
        RECT 273.745 95.860 274.170 96.320 ;
        RECT 270.465 95.430 271.315 95.680 ;
        RECT 266.810 95.225 268.465 95.430 ;
        RECT 266.810 95.080 267.040 95.225 ;
        RECT 205.335 91.970 207.495 93.150 ;
        RECT 252.335 92.800 254.495 93.980 ;
        RECT 262.635 92.460 262.895 95.080 ;
        RECT 263.155 94.850 263.575 95.030 ;
        RECT 266.185 94.850 266.605 95.030 ;
        RECT 263.155 94.800 266.615 94.850 ;
        RECT 263.175 94.645 266.615 94.800 ;
        RECT 267.715 93.915 267.935 95.225 ;
        RECT 268.175 95.175 268.465 95.225 ;
        RECT 267.715 93.820 270.865 93.915 ;
        RECT 267.715 93.695 270.895 93.820 ;
        RECT 267.715 92.865 267.935 93.695 ;
        RECT 270.475 93.590 270.895 93.695 ;
        RECT 271.080 93.755 273.595 94.005 ;
        RECT 270.085 93.405 270.315 93.540 ;
        RECT 266.165 92.645 267.935 92.865 ;
        RECT 268.215 93.200 270.315 93.405 ;
        RECT 266.185 92.510 266.605 92.645 ;
        RECT 205.335 90.310 207.495 91.490 ;
        RECT 252.335 91.140 254.495 92.320 ;
        RECT 262.635 92.000 262.950 92.460 ;
        RECT 266.810 92.310 267.040 92.460 ;
        RECT 268.215 92.310 268.420 93.200 ;
        RECT 270.085 93.080 270.315 93.200 ;
        RECT 270.475 92.935 270.895 93.030 ;
        RECT 271.080 92.935 271.330 93.755 ;
        RECT 273.165 93.590 273.585 93.755 ;
        RECT 273.880 93.540 274.170 95.860 ;
        RECT 274.480 93.935 274.675 101.680 ;
        RECT 283.225 100.575 285.385 101.760 ;
        RECT 330.225 101.320 332.385 102.500 ;
        RECT 283.255 100.540 285.360 100.575 ;
        RECT 283.225 98.920 285.385 100.105 ;
        RECT 330.225 99.660 332.385 100.840 ;
        RECT 283.255 98.880 285.360 98.920 ;
        RECT 283.225 97.265 285.385 98.450 ;
        RECT 330.225 98.000 332.385 99.180 ;
        RECT 283.255 97.220 285.360 97.265 ;
        RECT 283.225 95.610 285.385 96.795 ;
        RECT 330.225 96.340 332.385 97.520 ;
        RECT 283.255 95.560 285.360 95.610 ;
        RECT 283.225 93.955 285.385 95.140 ;
        RECT 330.225 94.680 332.385 95.860 ;
        RECT 274.480 93.740 277.230 93.935 ;
        RECT 283.255 93.900 285.360 93.955 ;
        RECT 276.795 93.580 277.215 93.740 ;
        RECT 273.745 93.080 274.170 93.540 ;
        RECT 277.455 93.530 277.735 93.570 ;
        RECT 270.460 92.685 271.330 92.935 ;
        RECT 266.810 92.105 268.420 92.310 ;
        RECT 266.810 92.000 267.040 92.105 ;
        RECT 205.335 88.650 207.495 89.830 ;
        RECT 252.335 89.480 254.495 90.660 ;
        RECT 262.635 89.380 262.895 92.000 ;
        RECT 263.155 91.720 263.575 91.950 ;
        RECT 266.185 91.720 266.605 91.950 ;
        RECT 263.175 91.515 266.615 91.720 ;
        RECT 267.740 91.145 267.960 92.105 ;
        RECT 267.740 90.925 270.915 91.145 ;
        RECT 271.080 90.935 273.595 91.185 ;
        RECT 267.740 89.865 267.960 90.925 ;
        RECT 270.475 90.810 270.895 90.925 ;
        RECT 270.475 90.140 270.895 90.250 ;
        RECT 271.080 90.140 271.330 90.935 ;
        RECT 273.165 90.810 273.585 90.935 ;
        RECT 273.880 90.760 274.170 93.080 ;
        RECT 277.375 93.070 277.735 93.530 ;
        RECT 273.745 90.300 274.170 90.760 ;
        RECT 277.455 90.750 277.735 93.070 ;
        RECT 283.225 92.300 285.385 93.485 ;
        RECT 330.225 93.020 332.385 94.200 ;
        RECT 283.255 92.240 285.360 92.300 ;
        RECT 270.475 90.020 271.330 90.140 ;
        RECT 270.480 89.890 271.330 90.020 ;
        RECT 266.170 89.645 267.960 89.865 ;
        RECT 266.185 89.430 266.605 89.645 ;
        RECT 262.635 89.140 262.950 89.380 ;
        RECT 205.335 86.990 207.495 88.170 ;
        RECT 252.335 87.820 254.495 89.000 ;
        RECT 262.630 88.920 262.950 89.140 ;
        RECT 262.630 88.890 262.895 88.920 ;
        RECT 205.335 85.330 207.495 86.510 ;
        RECT 252.335 86.160 254.495 87.340 ;
        RECT 262.630 87.280 262.890 88.890 ;
        RECT 263.155 88.725 263.575 88.870 ;
        RECT 266.185 88.725 266.605 88.870 ;
        RECT 263.155 88.640 266.605 88.725 ;
        RECT 263.160 88.520 266.600 88.640 ;
        RECT 269.265 88.260 270.855 88.485 ;
        RECT 269.265 88.225 270.895 88.260 ;
        RECT 269.265 87.280 269.525 88.225 ;
        RECT 270.475 88.030 270.895 88.225 ;
        RECT 271.080 88.215 273.605 88.465 ;
        RECT 273.880 88.380 274.170 90.300 ;
        RECT 277.375 90.290 277.735 90.750 ;
        RECT 283.225 90.645 285.385 91.830 ;
        RECT 330.225 91.360 332.385 92.540 ;
        RECT 283.255 90.580 285.360 90.645 ;
        RECT 273.880 88.250 277.190 88.380 ;
        RECT 262.630 87.020 269.525 87.280 ;
        RECT 269.990 87.520 270.315 87.980 ;
        RECT 263.255 86.580 263.495 87.020 ;
        RECT 266.290 86.580 266.535 87.020 ;
        RECT 263.155 86.350 263.575 86.580 ;
        RECT 266.185 86.350 266.605 86.580 ;
        RECT 266.900 86.300 267.160 87.020 ;
        RECT 262.720 86.290 262.950 86.300 ;
        RECT 262.655 85.840 262.950 86.290 ;
        RECT 266.810 85.840 267.160 86.300 ;
        RECT 252.335 84.500 254.495 85.680 ;
        RECT 262.655 84.085 262.865 85.840 ;
        RECT 266.900 85.815 267.160 85.840 ;
        RECT 269.990 86.540 270.260 87.520 ;
        RECT 270.475 87.405 270.895 87.470 ;
        RECT 271.080 87.405 271.330 88.215 ;
        RECT 273.165 88.030 273.585 88.215 ;
        RECT 273.880 88.160 277.215 88.250 ;
        RECT 273.880 87.980 274.170 88.160 ;
        RECT 276.795 88.020 277.215 88.160 ;
        RECT 273.745 87.520 274.170 87.980 ;
        RECT 277.455 87.970 277.735 90.290 ;
        RECT 283.225 88.990 285.385 90.175 ;
        RECT 330.225 89.700 332.385 90.880 ;
        RECT 283.255 88.920 285.360 88.990 ;
        RECT 270.475 87.240 271.330 87.405 ;
        RECT 270.500 87.155 271.330 87.240 ;
        RECT 269.990 86.155 270.975 86.540 ;
        RECT 269.990 85.200 270.260 86.155 ;
        RECT 273.880 85.680 274.170 87.520 ;
        RECT 277.375 87.510 277.735 87.970 ;
        RECT 277.455 86.115 277.735 87.510 ;
        RECT 283.225 87.335 285.385 88.520 ;
        RECT 330.225 88.040 332.385 89.220 ;
        RECT 283.255 87.260 285.360 87.335 ;
        RECT 277.455 86.020 278.375 86.115 ;
        RECT 277.455 85.740 278.410 86.020 ;
        RECT 270.470 85.590 274.170 85.680 ;
        RECT 277.490 85.660 278.375 85.740 ;
        RECT 283.225 85.680 285.385 86.865 ;
        RECT 330.225 86.380 332.385 87.560 ;
        RECT 283.255 85.600 285.360 85.680 ;
        RECT 270.470 85.470 277.170 85.590 ;
        RECT 270.470 85.395 277.215 85.470 ;
        RECT 270.475 85.250 270.895 85.395 ;
        RECT 273.165 85.250 273.585 85.395 ;
        RECT 273.880 85.315 277.215 85.395 ;
        RECT 273.880 85.200 274.170 85.315 ;
        RECT 276.795 85.240 277.215 85.315 ;
        RECT 269.990 84.740 270.315 85.200 ;
        RECT 273.745 84.815 274.170 85.200 ;
        RECT 273.745 84.740 273.975 84.815 ;
        RECT 262.025 83.745 263.010 84.085 ;
        RECT 265.955 83.735 267.315 83.830 ;
        RECT 269.990 83.735 270.260 84.740 ;
        RECT 270.475 84.460 270.895 84.690 ;
        RECT 275.310 84.555 275.650 85.140 ;
        RECT 277.375 85.090 277.605 85.190 ;
        RECT 278.610 85.090 278.950 85.140 ;
        RECT 277.375 84.830 278.950 85.090 ;
        RECT 277.375 84.730 277.605 84.830 ;
        RECT 276.795 84.555 277.215 84.680 ;
        RECT 265.955 83.465 270.260 83.735 ;
        RECT 270.530 83.765 270.830 84.460 ;
        RECT 275.310 84.450 277.215 84.555 ;
        RECT 275.310 84.305 277.195 84.450 ;
        RECT 275.310 84.050 275.650 84.305 ;
        RECT 278.610 84.040 278.950 84.830 ;
        RECT 283.225 84.025 285.385 85.210 ;
        RECT 330.225 84.720 332.385 85.900 ;
        RECT 283.255 83.940 285.360 84.025 ;
        RECT 270.530 83.465 282.235 83.765 ;
        RECT 265.955 83.355 267.315 83.465 ;
        RECT 275.275 83.190 276.220 83.265 ;
        RECT 270.520 83.090 276.220 83.190 ;
        RECT 277.270 83.125 278.155 83.215 ;
        RECT 264.865 82.865 276.220 83.090 ;
        RECT 264.865 82.765 270.790 82.865 ;
        RECT 275.275 82.810 276.220 82.865 ;
        RECT 276.690 82.825 278.155 83.125 ;
        RECT 264.865 82.740 265.220 82.765 ;
        RECT 258.525 82.440 265.220 82.740 ;
        RECT 276.690 82.625 276.990 82.825 ;
        RECT 277.270 82.760 278.155 82.825 ;
        RECT 254.115 82.415 265.220 82.440 ;
        RECT 254.115 82.115 259.105 82.415 ;
        RECT 271.050 82.325 276.990 82.625 ;
        RECT 262.220 82.120 263.105 82.205 ;
        RECT 205.385 80.670 207.545 81.850 ;
        RECT 254.115 81.800 254.440 82.115 ;
        RECT 252.410 81.550 254.515 81.800 ;
        RECT 262.220 81.765 263.110 82.120 ;
        RECT 271.050 82.105 271.350 82.325 ;
        RECT 205.385 79.010 207.545 80.190 ;
        RECT 252.385 79.840 254.545 81.020 ;
        RECT 261.160 80.520 262.160 81.520 ;
        RECT 205.385 77.350 207.545 78.530 ;
        RECT 252.385 78.180 254.545 79.360 ;
        RECT 261.470 79.100 261.710 80.520 ;
        RECT 262.805 80.260 263.110 81.765 ;
        RECT 264.495 81.795 271.350 82.105 ;
        RECT 278.625 82.080 278.965 82.990 ;
        RECT 272.105 81.890 278.965 82.080 ;
        RECT 264.495 81.520 264.805 81.795 ;
        RECT 272.105 81.780 278.960 81.890 ;
        RECT 263.850 80.520 264.850 81.520 ;
        RECT 272.105 81.490 272.405 81.780 ;
        RECT 262.220 79.955 263.110 80.260 ;
        RECT 259.320 78.880 259.550 79.010 ;
        RECT 260.290 78.880 260.520 79.010 ;
        RECT 261.430 78.880 261.760 79.100 ;
        RECT 259.320 78.680 261.760 78.880 ;
        RECT 259.320 78.550 259.550 78.680 ;
        RECT 260.290 78.550 260.520 78.680 ;
        RECT 261.430 78.510 261.760 78.680 ;
        RECT 259.710 78.310 260.130 78.500 ;
        RECT 262.220 78.310 262.525 79.955 ;
        RECT 264.480 79.790 264.810 80.520 ;
        RECT 265.590 80.490 266.590 81.490 ;
        RECT 271.450 80.490 272.450 81.490 ;
        RECT 273.190 80.520 274.190 81.520 ;
        RECT 275.880 80.520 276.880 81.520 ;
        RECT 265.630 79.790 265.960 80.490 ;
        RECT 272.080 79.790 272.410 80.490 ;
        RECT 273.230 79.790 273.560 80.520 ;
        RECT 263.210 79.300 266.970 79.590 ;
        RECT 271.070 79.300 274.830 79.590 ;
        RECT 263.205 79.260 266.975 79.300 ;
        RECT 262.720 78.860 263.050 79.090 ;
        RECT 263.205 79.070 263.625 79.260 ;
        RECT 266.555 79.070 266.975 79.260 ;
        RECT 271.065 79.260 274.835 79.300 ;
        RECT 271.065 79.070 271.485 79.260 ;
        RECT 274.415 79.070 274.835 79.260 ;
        RECT 276.330 79.100 276.570 80.520 ;
        RECT 263.830 78.860 264.060 79.020 ;
        RECT 266.120 78.930 266.350 79.020 ;
        RECT 267.180 78.930 267.410 79.020 ;
        RECT 262.720 78.650 264.140 78.860 ;
        RECT 265.620 78.670 267.410 78.930 ;
        RECT 262.720 78.500 263.050 78.650 ;
        RECT 263.830 78.560 264.060 78.650 ;
        RECT 263.205 78.310 263.625 78.510 ;
        RECT 265.620 78.380 265.880 78.670 ;
        RECT 266.120 78.560 266.350 78.670 ;
        RECT 267.180 78.560 267.410 78.670 ;
        RECT 270.630 78.930 270.860 79.020 ;
        RECT 271.690 78.930 271.920 79.020 ;
        RECT 270.630 78.670 272.420 78.930 ;
        RECT 273.980 78.860 274.210 79.020 ;
        RECT 274.990 78.860 275.320 79.090 ;
        RECT 270.630 78.560 270.860 78.670 ;
        RECT 271.690 78.560 271.920 78.670 ;
        RECT 272.160 78.380 272.420 78.670 ;
        RECT 273.900 78.650 275.320 78.860 ;
        RECT 273.980 78.560 274.210 78.650 ;
        RECT 263.810 78.310 264.140 78.380 ;
        RECT 265.590 78.310 265.920 78.380 ;
        RECT 259.670 78.050 265.920 78.310 ;
        RECT 263.810 77.790 264.140 78.050 ;
        RECT 265.590 77.790 265.920 78.050 ;
        RECT 272.120 78.310 272.450 78.380 ;
        RECT 273.900 78.310 274.230 78.380 ;
        RECT 274.415 78.310 274.835 78.510 ;
        RECT 274.990 78.500 275.320 78.650 ;
        RECT 276.280 78.880 276.610 79.100 ;
        RECT 277.520 78.880 277.750 79.010 ;
        RECT 278.490 78.880 278.720 79.010 ;
        RECT 276.280 78.680 278.720 78.880 ;
        RECT 276.280 78.510 276.610 78.680 ;
        RECT 277.520 78.550 277.750 78.680 ;
        RECT 278.490 78.550 278.720 78.680 ;
        RECT 277.910 78.310 278.330 78.500 ;
        RECT 272.120 78.050 278.370 78.310 ;
        RECT 272.120 77.790 272.450 78.050 ;
        RECT 273.900 77.790 274.230 78.050 ;
        RECT 205.385 75.690 207.545 76.870 ;
        RECT 252.385 76.520 254.545 77.700 ;
        RECT 262.720 76.460 263.050 76.740 ;
        RECT 264.470 76.460 264.800 76.730 ;
        RECT 273.240 76.460 273.570 76.730 ;
        RECT 274.990 76.460 275.320 76.740 ;
        RECT 259.690 76.200 265.890 76.460 ;
        RECT 205.385 74.030 207.545 75.210 ;
        RECT 252.385 74.860 254.545 76.040 ;
        RECT 259.700 76.030 260.120 76.200 ;
        RECT 262.720 76.150 263.050 76.200 ;
        RECT 263.215 76.020 263.635 76.200 ;
        RECT 264.470 76.140 264.800 76.200 ;
        RECT 262.780 75.860 263.010 75.970 ;
        RECT 263.820 75.860 264.150 76.040 ;
        RECT 262.780 75.650 264.150 75.860 ;
        RECT 262.780 75.510 263.010 75.650 ;
        RECT 263.215 75.250 263.635 75.460 ;
        RECT 263.820 75.450 264.150 75.650 ;
        RECT 265.630 75.840 265.890 76.200 ;
        RECT 272.150 76.200 278.350 76.460 ;
        RECT 266.120 75.840 266.350 75.940 ;
        RECT 267.180 75.840 267.410 75.940 ;
        RECT 265.630 75.580 267.410 75.840 ;
        RECT 266.120 75.480 266.350 75.580 ;
        RECT 267.180 75.480 267.410 75.580 ;
        RECT 270.630 75.840 270.860 75.940 ;
        RECT 271.690 75.840 271.920 75.940 ;
        RECT 272.150 75.840 272.410 76.200 ;
        RECT 273.240 76.140 273.570 76.200 ;
        RECT 270.630 75.580 272.410 75.840 ;
        RECT 273.890 75.860 274.220 76.040 ;
        RECT 274.405 76.020 274.825 76.200 ;
        RECT 274.990 76.150 275.320 76.200 ;
        RECT 277.920 76.030 278.340 76.200 ;
        RECT 275.030 75.860 275.260 75.970 ;
        RECT 273.890 75.650 275.260 75.860 ;
        RECT 270.630 75.480 270.860 75.580 ;
        RECT 271.690 75.480 271.920 75.580 ;
        RECT 273.890 75.450 274.220 75.650 ;
        RECT 275.030 75.510 275.260 75.650 ;
        RECT 266.555 75.250 266.975 75.430 ;
        RECT 263.210 75.200 266.975 75.250 ;
        RECT 271.065 75.250 271.485 75.430 ;
        RECT 274.405 75.250 274.825 75.460 ;
        RECT 271.065 75.200 274.830 75.250 ;
        RECT 263.210 74.920 266.970 75.200 ;
        RECT 271.070 74.920 274.830 75.200 ;
        RECT 205.385 72.370 207.545 73.550 ;
        RECT 252.385 73.200 254.545 74.380 ;
        RECT 205.385 70.710 207.545 71.890 ;
        RECT 252.385 71.540 254.545 72.720 ;
        RECT 205.385 69.050 207.545 70.230 ;
        RECT 252.385 69.880 254.545 71.060 ;
        RECT 274.050 70.920 276.155 70.960 ;
        RECT 274.050 70.430 280.035 70.920 ;
        RECT 274.050 70.370 276.155 70.430 ;
        RECT 205.385 67.390 207.545 68.570 ;
        RECT 252.385 68.220 254.545 69.400 ;
        RECT 261.430 67.970 261.760 68.460 ;
        RECT 267.845 68.110 268.105 68.660 ;
        RECT 261.400 67.810 265.250 67.970 ;
        RECT 261.030 67.760 265.250 67.810 ;
        RECT 252.385 66.560 254.545 67.740 ;
        RECT 261.030 67.580 262.030 67.760 ;
        RECT 264.220 67.580 265.220 67.760 ;
        RECT 267.850 67.195 268.050 68.110 ;
        RECT 276.280 67.970 276.610 68.460 ;
        RECT 272.790 67.810 276.640 67.970 ;
        RECT 272.790 67.760 277.010 67.810 ;
        RECT 272.820 67.580 273.820 67.760 ;
        RECT 276.010 67.580 277.010 67.760 ;
        RECT 267.850 67.160 268.085 67.195 ;
        RECT 266.950 66.950 268.085 67.160 ;
        RECT 265.110 65.075 265.340 65.130 ;
        RECT 266.950 65.075 267.150 66.950 ;
        RECT 267.855 66.905 268.085 66.950 ;
        RECT 268.245 66.715 268.745 66.945 ;
        RECT 268.340 65.320 268.565 66.715 ;
        RECT 270.125 66.405 270.400 66.775 ;
        RECT 268.245 65.090 268.745 65.320 ;
        RECT 270.175 65.130 270.345 66.405 ;
        RECT 279.545 65.765 280.035 70.430 ;
        RECT 281.935 66.810 282.235 83.465 ;
        RECT 283.225 82.370 285.385 83.555 ;
        RECT 330.225 83.060 332.385 84.240 ;
        RECT 283.255 82.280 285.360 82.370 ;
        RECT 283.225 80.715 285.385 81.900 ;
        RECT 330.225 81.400 332.385 82.580 ;
        RECT 283.255 80.620 285.360 80.715 ;
        RECT 283.225 79.060 285.385 80.245 ;
        RECT 330.225 79.740 332.385 80.920 ;
        RECT 283.255 78.960 285.360 79.060 ;
        RECT 283.225 77.405 285.385 78.590 ;
        RECT 330.225 78.080 332.385 79.260 ;
        RECT 283.255 77.300 285.360 77.405 ;
        RECT 283.225 75.750 285.385 76.935 ;
        RECT 330.225 76.420 332.385 77.600 ;
        RECT 283.255 75.640 285.360 75.750 ;
        RECT 283.225 74.095 285.385 75.280 ;
        RECT 330.225 74.760 332.385 75.940 ;
        RECT 283.255 73.980 285.360 74.095 ;
        RECT 283.225 72.440 285.385 73.625 ;
        RECT 330.225 73.100 332.385 74.280 ;
        RECT 283.255 72.320 285.360 72.440 ;
        RECT 283.225 70.785 285.385 71.970 ;
        RECT 330.225 71.440 332.385 72.620 ;
        RECT 283.255 70.660 285.360 70.785 ;
        RECT 283.225 69.130 285.385 70.315 ;
        RECT 330.225 69.780 332.385 70.960 ;
        RECT 283.255 69.000 285.360 69.130 ;
        RECT 283.225 67.475 285.385 68.660 ;
        RECT 330.225 68.120 332.385 69.300 ;
        RECT 283.255 67.340 285.360 67.475 ;
        RECT 281.935 66.460 285.385 66.810 ;
        RECT 330.225 66.460 332.385 67.640 ;
        RECT 271.155 65.275 280.035 65.765 ;
        RECT 263.905 64.690 264.905 64.880 ;
        RECT 265.110 64.875 267.150 65.075 ;
        RECT 265.110 64.840 265.340 64.875 ;
        RECT 268.245 64.690 268.745 64.880 ;
        RECT 270.145 64.840 270.375 65.130 ;
        RECT 270.535 64.690 270.955 64.880 ;
        RECT 271.155 64.690 271.645 65.275 ;
        RECT 263.890 64.195 271.645 64.690 ;
      LAYER via ;
        RECT 268.770 100.545 269.030 100.805 ;
        RECT 269.090 100.545 269.350 100.805 ;
        RECT 267.225 99.300 267.485 99.560 ;
        RECT 267.545 99.300 267.805 99.560 ;
        RECT 267.865 99.300 268.125 99.560 ;
        RECT 268.310 98.670 268.570 98.930 ;
        RECT 268.630 98.670 268.890 98.930 ;
        RECT 270.310 97.375 270.570 97.635 ;
        RECT 270.630 97.375 270.890 97.635 ;
        RECT 268.190 95.880 268.450 96.140 ;
        RECT 268.190 95.560 268.450 95.820 ;
        RECT 268.190 95.240 268.450 95.500 ;
        RECT 270.270 86.220 270.530 86.480 ;
        RECT 270.590 86.220 270.850 86.480 ;
        RECT 277.645 85.760 277.905 86.020 ;
        RECT 277.965 85.760 278.225 86.020 ;
        RECT 275.350 84.790 275.610 85.050 ;
        RECT 262.230 83.785 262.490 84.045 ;
        RECT 262.550 83.785 262.810 84.045 ;
        RECT 278.650 84.780 278.910 85.040 ;
        RECT 275.350 84.470 275.610 84.730 ;
        RECT 266.025 83.465 266.285 83.725 ;
        RECT 266.345 83.465 266.605 83.725 ;
        RECT 266.665 83.465 266.925 83.725 ;
        RECT 266.985 83.465 267.245 83.725 ;
        RECT 278.650 84.460 278.910 84.720 ;
        RECT 275.350 84.150 275.610 84.410 ;
        RECT 278.650 84.140 278.910 84.400 ;
        RECT 275.490 82.910 275.750 83.170 ;
        RECT 275.810 82.910 276.070 83.170 ;
        RECT 277.425 82.860 277.685 83.120 ;
        RECT 277.745 82.860 278.005 83.120 ;
        RECT 278.665 82.630 278.925 82.890 ;
        RECT 262.375 81.855 262.635 82.115 ;
        RECT 262.695 81.855 262.955 82.115 ;
        RECT 278.665 82.310 278.925 82.570 ;
        RECT 278.665 81.990 278.925 82.250 ;
        RECT 264.515 79.955 264.775 80.215 ;
        RECT 261.465 78.675 261.725 78.935 ;
        RECT 265.665 79.955 265.925 80.215 ;
        RECT 272.115 79.955 272.375 80.215 ;
        RECT 273.265 79.955 273.525 80.215 ;
        RECT 262.755 78.665 263.015 78.925 ;
        RECT 275.025 78.665 275.285 78.925 ;
        RECT 263.845 77.955 264.105 78.215 ;
        RECT 265.625 77.955 265.885 78.215 ;
        RECT 276.315 78.675 276.575 78.935 ;
        RECT 272.155 77.955 272.415 78.215 ;
        RECT 273.935 77.955 274.195 78.215 ;
        RECT 262.755 76.315 263.015 76.575 ;
        RECT 264.505 76.305 264.765 76.565 ;
        RECT 263.855 75.615 264.115 75.875 ;
        RECT 273.275 76.305 273.535 76.565 ;
        RECT 275.025 76.315 275.285 76.575 ;
        RECT 273.925 75.615 274.185 75.875 ;
        RECT 261.465 68.035 261.725 68.295 ;
        RECT 267.845 68.255 268.105 68.515 ;
        RECT 276.315 68.035 276.575 68.295 ;
        RECT 270.135 66.460 270.395 66.720 ;
      LAYER met2 ;
        RECT 268.615 100.525 269.505 100.820 ;
        RECT 267.165 99.265 268.185 99.590 ;
        RECT 267.540 85.080 267.800 99.265 ;
        RECT 268.685 98.945 268.910 100.525 ;
        RECT 268.155 98.650 269.045 98.945 ;
        RECT 268.215 96.155 268.440 98.650 ;
        RECT 270.130 97.360 271.065 97.645 ;
        RECT 268.125 95.225 268.515 96.155 ;
        RECT 270.225 86.490 270.530 97.360 ;
        RECT 270.090 86.205 271.025 86.490 ;
        RECT 277.440 85.710 278.425 86.065 ;
        RECT 267.540 84.820 268.510 85.080 ;
        RECT 262.075 83.780 263.010 84.135 ;
        RECT 262.075 83.695 267.365 83.780 ;
        RECT 262.560 83.410 267.365 83.695 ;
        RECT 262.560 82.155 262.995 83.410 ;
        RECT 265.925 83.405 267.365 83.410 ;
        RECT 262.170 81.815 263.155 82.155 ;
        RECT 264.430 79.840 264.860 80.330 ;
        RECT 265.580 79.840 266.010 80.330 ;
        RECT 261.380 78.560 261.810 79.050 ;
        RECT 261.460 69.000 261.730 78.560 ;
        RECT 262.670 78.550 263.100 79.040 ;
        RECT 262.770 76.690 263.040 78.550 ;
        RECT 263.840 78.330 264.110 78.400 ;
        RECT 263.760 77.840 264.190 78.330 ;
        RECT 262.670 76.200 263.100 76.690 ;
        RECT 262.770 76.100 263.040 76.200 ;
        RECT 263.840 75.990 264.110 77.840 ;
        RECT 264.490 76.680 264.770 79.840 ;
        RECT 265.650 78.330 265.920 79.840 ;
        RECT 265.540 77.840 265.970 78.330 ;
        RECT 264.420 76.190 264.850 76.680 ;
        RECT 263.770 75.500 264.200 75.990 ;
        RECT 268.250 72.155 268.510 84.820 ;
        RECT 275.260 84.100 275.700 85.100 ;
        RECT 275.285 83.215 275.650 84.100 ;
        RECT 275.275 82.860 276.275 83.215 ;
        RECT 277.625 83.165 277.935 85.710 ;
        RECT 278.560 84.090 279.000 85.090 ;
        RECT 277.220 82.810 278.205 83.165 ;
        RECT 278.645 82.940 278.935 84.090 ;
        RECT 278.575 81.940 279.015 82.940 ;
        RECT 272.030 79.840 272.460 80.330 ;
        RECT 273.180 79.840 273.610 80.330 ;
        RECT 272.120 78.330 272.390 79.840 ;
        RECT 272.070 77.840 272.500 78.330 ;
        RECT 273.270 76.680 273.550 79.840 ;
        RECT 274.940 78.550 275.370 79.040 ;
        RECT 276.230 78.560 276.660 79.050 ;
        RECT 273.930 78.330 274.200 78.400 ;
        RECT 273.850 77.840 274.280 78.330 ;
        RECT 273.190 76.190 273.620 76.680 ;
        RECT 273.930 75.990 274.200 77.840 ;
        RECT 275.000 76.690 275.270 78.550 ;
        RECT 274.940 76.200 275.370 76.690 ;
        RECT 275.000 76.100 275.270 76.200 ;
        RECT 273.840 75.500 274.270 75.990 ;
        RECT 267.850 71.895 268.510 72.155 ;
        RECT 261.460 68.410 261.775 69.000 ;
        RECT 267.850 68.610 268.110 71.895 ;
        RECT 261.380 67.920 261.810 68.410 ;
        RECT 267.795 68.160 268.150 68.610 ;
        RECT 276.310 68.410 276.580 78.560 ;
        RECT 276.230 67.920 276.660 68.410 ;
        RECT 261.505 66.725 261.775 67.920 ;
        RECT 261.505 66.455 270.465 66.725 ;
  END
END sky130_ef_ip__xtal_osc_32k_DI
END LIBRARY

